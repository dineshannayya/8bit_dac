* C:\FOSSEE\eSim\library\SubcircuitLibrary\2bit_DAC\2bit_DAC.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 04/22/23 17:36:35

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
U1  /vdd /d0 /d1 /vrefh /vrefl /vout Net-_S1-Pad7_ PORT		
R1  /vrefh Net-_R1-Pad2_ resistor		
S1  /vdd /d0 /vrefl Net-_R1-Pad2_ Net-_S1-Pad5_ Net-_S1-Pad6_ Net-_S1-Pad7_ switch_2n		
S2  /vdd /d1 Net-_S1-Pad6_ Net-_S1-Pad5_ /vout switch		

.end
