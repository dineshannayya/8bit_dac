* SPICE3 file created from switch.ext - technology: sky130B

.lib "sky130_fd_pr/models/sky130.lib.spice" tt


.subckt switch vrefh vrefl Vout D1 vdd gnd
X0 a_n310_n202# D1 gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.116e+11p ps=3.64e+06u w=420000u l=500000u
X1 Vout a_n310_n202# vrefl gnd sky130_fd_pr__nfet_01v8 ad=3.696e+11p pd=3.44e+06u as=2.058e+11p ps=1.82e+06u w=420000u l=500000u
X2 a_116_n202# a_n310_n202# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=500000u
X3 vrefh a_116_n202# Vout gnd sky130_fd_pr__nfet_01v8 ad=2.058e+11p pd=1.82e+06u as=0p ps=0u w=420000u l=500000u
X4 a_n310_n202# D1 vdd vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=8.8e+11p ps=5.76e+06u w=1e+06u l=500000u
X5 a_116_n202# a_n310_n202# vdd vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X6 vrefl a_116_n202# Vout vdd sky130_fd_pr__pfet_01v8 ad=4.431e+11p pd=2.9e+06u as=8.4e+11p ps=5.68e+06u w=1e+06u l=500000u
X7 Vout a_n310_n202# vrefh vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=4.4e+11p ps=2.88e+06u w=1e+06u l=500000u
C0 vdd gnd 3.36fF
.ends

Xsub1 vrefh vrefl Vout D1 vdd gnd switch

Vdd vdd 0 dc 1.8
Vin1 vrefh 0 dc 2.5
Vin2 vrefl 0 dc 2.2
Vd0 D1 0 pulse(0 1.8 0ns 0.1ns 0.1ns 5ns 10ns)

.tran 0.1ns 20ns
.control
run
plot V(vout) V(D1)
.endc
.end
