* D:\vlsi\github\8bit_dac\schematics\2bit_DAC\2bit_DAC.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 04/19/23 16:29:56

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
R4  Net-_R3-Pad2_ /vrefl resistor		
R3  Net-_R2-Pad2_ Net-_R3-Pad2_ resistor		
R2  Net-_R1-Pad2_ Net-_R2-Pad2_ resistor		
R1  /vrefh Net-_R1-Pad2_ resistor		
U1  /vdd /vrefh /vrefl /d0 /d1 /vout PORT		
S2  /vdd /d0 Net-_R3-Pad2_ /vrefl Net-_S2-Pad5_ switch		
S1  /vdd /d0 Net-_R1-Pad2_ Net-_R2-Pad2_ Net-_S1-Pad5_ switch		
S3  /vdd /d1 Net-_S1-Pad5_ Net-_S2-Pad5_ /vout switch		

.end
