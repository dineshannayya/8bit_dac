* SPICE3 file created from switch2n.ext - technology: sky130B

.lib "sky130_fd_pr/models/sky130.lib.spice" tt

.subckt switch2n vrefh0 vrefl0 vrefh1 D0_INV vrefl1 D0_BUF Vout0 Vout1 D0 vdd gnd
X0 vrefh0 D0_BUF Vout0 gnd sky130_fd_pr__nfet_01v8 ad=2.058e+11p pd=1.82e+06u as=3.696e+11p ps=3.44e+06u w=420000u l=500000u
X1 D0_BUF D0_INV vdd vdd sky130_fd_pr__pfet_01v8 ad=4.2e+11p pd=2.84e+06u as=8.8e+11p ps=5.76e+06u w=1e+06u l=500000u
X2 Vout1 D0_INV vrefl1 gnd sky130_fd_pr__nfet_01v8 ad=3.696e+11p pd=3.44e+06u as=2.058e+11p ps=1.82e+06u w=420000u l=500000u
X3 D0_INV D0 vdd vdd sky130_fd_pr__pfet_01v8 ad=4.2e+11p pd=2.84e+06u as=0p ps=0u w=1e+06u l=500000u
X4 D0_BUF D0_INV gnd gnd sky130_fd_pr__nfet_01v8 ad=1.848e+11p pd=1.72e+06u as=4.116e+11p ps=3.64e+06u w=420000u l=500000u
X5 D0_INV D0 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.848e+11p pd=1.72e+06u as=0p ps=0u w=420000u l=500000u
X6 vrefl0 D0_BUF Vout0 vdd sky130_fd_pr__pfet_01v8 ad=4.431e+11p pd=2.9e+06u as=8.4e+11p ps=5.68e+06u w=1e+06u l=500000u
X7 Vout0 D0_INV vrefh0 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=4.4e+11p ps=2.88e+06u w=1e+06u l=500000u
X8 Vout1 D0_INV vrefh1 vdd sky130_fd_pr__pfet_01v8 ad=8.4e+11p pd=5.68e+06u as=4.4e+11p ps=2.88e+06u w=1e+06u l=500000u
X9 vrefh1 D0_BUF Vout1 gnd sky130_fd_pr__nfet_01v8 ad=2.058e+11p pd=1.82e+06u as=0p ps=0u w=420000u l=500000u
X10 Vout0 D0_INV vrefl0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.058e+11p ps=1.82e+06u w=420000u l=500000u
X11 vrefl1 D0_BUF Vout1 vdd sky130_fd_pr__pfet_01v8 ad=4.431e+11p pd=2.9e+06u as=0p ps=0u w=1e+06u l=500000u
C0 vdd gnd 4.61fF
.ends
Xsub1 vrefh0 vrefl0 vrefh1 D0_INV vrefl1 D0_BUF Vout0 Vout1 D0 vdd gnd switch2n

Vdd vdd 0 dc 1.8
Vin1 vrefh0 0 dc 2.5
Vin2 vrefl0 0 dc 2.2
Vin3 vrefh1 0 dc 1.5
Vin4 vrefl1 0 dc 1.2
Vd0 D0 0 pulse(0 1.8 0ns 0.1ns 0.1ns 5ns 10ns)

.tran 0.1ns 20ns
.control
run
plot V(Vout0) V(Vout1) V(D0) 
* plot V(D0) V(D0_INV) V(D0_BUF)
.endc
.end



