module dac_top (Vout0,
    Vout1,
    Vout2,
    Vout3,
    Vref,
    vdda1,
    vssa1,
    DIn0,
    DIn1,
    DIn2,
    DIn3);
 output Vout0;
 output Vout1;
 output Vout2;
 output Vout3;
 input Vref;
 input vdda1;
 input vssa1;
 input [7:0] DIn0;
 input [7:0] DIn1;
 input [7:0] DIn2;
 input [7:0] DIn3;

 wire clknet_0_Vref;
 wire clknet_1_0__leaf_Vref;
 wire clknet_1_1__leaf_Vref;

 sky130_fd_sc_hd__diode_2 ANTENNA__0__CLK (.DIODE(clknet_1_1__leaf_Vref),
    .VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__diode_2 ANTENNA__0__D (.DIODE(DIn1[7]),
    .VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__diode_2 ANTENNA__1__CLK (.DIODE(clknet_1_1__leaf_Vref),
    .VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__diode_2 ANTENNA__1__D (.DIODE(DIn2[7]),
    .VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__diode_2 ANTENNA__2__CLK (.DIODE(clknet_1_0__leaf_Vref),
    .VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__diode_2 ANTENNA__2__D (.DIODE(DIn0[0]),
    .VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__diode_2 ANTENNA__3__CLK (.DIODE(clknet_1_0__leaf_Vref),
    .VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__diode_2 ANTENNA__3__D (.DIODE(DIn1[0]),
    .VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_Vref_A (.DIODE(Vref),
    .VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_Vref_A (.DIODE(clknet_0_Vref),
    .VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_Vref_A (.DIODE(clknet_0_Vref),
    .VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_0_109 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_0_113 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_0_125 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_0_137 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_0_141 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_0_15 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_0_153 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_0_165 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_0_169 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_0_181 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_0_193 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_0_197 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_0_209 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_0_221 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_0_225 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_0_237 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_0_249 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_0_253 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_0_265 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_0_27 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_0_277 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_0_281 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_0_29 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_0_293 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_0_3 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_0_305 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_0_309 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_0_321 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_0_333 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_0_337 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_0_349 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_0_361 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_0_365 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_0_377 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_0_389 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_0_393 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_0_405 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_0_41 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_0_417 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_0_421 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_0_433 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_0_445 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_0_449 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_0_461 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_0_473 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_0_477 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_0_489 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_0_501 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_8 FILLER_0_505 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_0_513 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_0_53 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_0_57 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_0_69 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_0_81 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_0_85 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_0_97 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_100_109 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_100_121 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_100_133 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_100_139 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_100_141 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_100_15 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_100_153 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_100_165 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_100_177 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_100_189 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_100_195 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_100_197 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_100_209 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_100_221 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_100_233 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_100_245 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_100_251 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_100_253 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_100_265 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_100_27 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_100_277 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_100_289 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_100_29 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_100_3 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_100_301 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_100_307 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_100_309 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_100_321 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_100_333 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_100_345 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_100_357 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_100_363 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_100_365 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_100_377 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_100_389 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_100_401 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_100_41 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_100_413 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_100_419 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_100_421 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_100_433 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_100_445 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_100_457 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_100_469 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_100_475 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_100_477 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_100_489 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_100_501 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_100_513 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_100_53 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_100_65 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_100_77 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_100_83 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_100_85 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_100_97 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_101_105 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_101_111 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_101_113 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_101_125 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_101_137 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_101_149 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_101_15 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_101_161 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_101_167 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_101_169 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_101_181 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_101_193 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_101_205 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_101_217 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_101_223 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_101_225 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_101_237 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_101_249 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_101_261 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_101_27 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_101_273 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_101_279 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_101_281 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_101_293 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_101_3 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_101_305 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_101_317 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_101_329 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_101_335 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_101_337 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_101_349 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_101_361 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_101_373 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_101_385 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_101_39 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_101_391 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_101_393 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_101_405 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_101_417 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_101_429 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_101_441 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_101_447 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_101_449 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_101_461 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_101_473 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_101_485 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_101_497 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_101_503 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_8 FILLER_101_505 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_4 FILLER_101_51 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_101_513 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_101_55 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_101_57 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_101_69 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_101_81 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_101_93 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_102_109 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_102_121 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_102_133 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_102_139 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_102_141 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_102_15 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_102_153 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_102_165 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_102_177 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_102_189 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_102_195 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_102_197 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_102_209 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_102_221 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_102_233 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_102_245 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_102_251 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_102_253 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_102_265 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_102_27 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_102_277 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_102_289 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_102_29 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_102_3 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_102_301 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_102_307 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_102_309 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_102_321 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_102_333 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_102_345 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_102_357 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_102_363 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_102_365 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_102_377 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_102_389 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_102_401 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_102_41 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_102_413 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_102_419 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_102_421 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_102_433 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_102_445 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_102_457 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_102_469 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_102_475 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_102_477 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_102_489 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_102_501 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_102_513 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_102_53 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_102_65 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_102_77 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_102_83 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_102_85 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_102_97 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_103_105 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_103_111 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_103_113 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_103_125 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_103_137 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_103_149 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_103_15 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_103_161 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_103_167 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_103_169 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_103_181 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_103_193 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_103_205 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_103_217 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_103_223 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_103_225 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_103_237 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_103_249 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_103_261 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_103_27 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_103_273 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_103_279 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_103_281 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_103_293 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_103_3 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_103_305 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_103_317 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_103_329 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_103_335 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_103_337 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_103_349 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_103_361 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_103_373 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_103_385 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_103_39 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_103_391 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_103_393 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_103_405 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_103_417 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_103_429 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_103_441 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_103_447 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_103_449 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_103_461 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_103_473 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_103_485 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_103_497 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_103_503 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_8 FILLER_103_505 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_4 FILLER_103_51 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_103_513 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_103_55 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_103_57 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_103_69 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_103_81 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_103_93 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_104_109 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_104_121 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_104_133 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_104_139 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_104_141 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_104_15 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_104_153 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_104_165 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_104_177 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_104_189 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_104_195 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_104_197 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_104_209 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_104_221 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_104_233 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_104_245 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_104_251 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_104_253 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_104_265 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_104_27 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_104_277 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_104_289 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_104_29 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_104_3 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_104_301 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_104_307 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_104_309 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_104_321 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_104_333 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_104_345 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_104_357 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_104_363 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_104_365 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_104_377 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_104_389 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_104_401 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_104_41 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_104_413 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_104_419 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_104_421 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_104_433 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_104_445 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_104_457 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_104_469 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_104_475 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_104_477 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_104_489 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_104_501 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_104_513 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_104_53 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_104_65 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_104_77 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_104_83 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_104_85 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_104_97 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_105_105 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_105_111 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_105_113 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_105_125 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_105_137 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_105_149 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_105_15 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_105_161 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_105_167 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_105_169 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_105_181 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_105_193 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_105_205 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_105_217 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_105_223 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_105_225 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_105_237 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_105_249 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_105_261 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_105_27 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_105_273 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_105_279 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_105_281 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_105_293 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_105_3 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_105_305 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_105_317 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_105_329 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_105_335 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_105_337 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_105_349 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_105_361 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_105_373 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_105_385 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_105_39 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_105_391 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_105_393 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_105_405 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_105_417 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_105_429 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_105_441 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_105_447 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_105_449 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_105_461 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_105_473 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_105_485 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_105_497 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_105_503 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_8 FILLER_105_505 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_4 FILLER_105_51 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_105_513 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_105_55 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_105_57 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_105_69 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_105_81 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_105_93 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_106_109 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_106_121 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_106_133 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_106_139 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_106_141 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_106_15 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_106_153 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_106_165 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_106_177 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_106_189 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_106_195 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_106_197 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_106_209 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_106_221 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_106_233 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_106_245 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_106_251 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_106_253 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_106_265 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_106_27 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_106_277 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_106_289 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_106_29 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_106_3 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_106_301 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_106_307 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_106_309 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_106_321 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_106_333 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_106_345 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_106_357 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_106_363 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_106_365 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_106_377 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_106_389 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_106_401 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_106_41 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_106_413 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_106_419 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_106_421 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_106_433 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_106_445 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_106_457 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_106_469 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_106_475 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_106_477 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_106_489 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_106_501 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_106_513 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_106_53 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_106_65 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_106_77 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_106_83 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_106_85 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_106_97 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_107_105 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_107_111 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_107_113 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_107_125 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_107_137 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_107_149 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_107_15 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_107_161 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_107_167 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_107_169 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_107_181 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_107_193 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_107_205 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_107_217 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_107_223 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_107_225 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_107_237 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_107_249 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_107_261 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_107_27 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_107_273 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_107_279 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_107_281 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_107_293 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_107_3 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_107_305 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_107_317 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_107_329 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_107_335 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_107_337 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_107_349 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_107_361 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_107_373 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_107_385 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_107_39 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_107_391 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_107_393 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_107_405 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_107_417 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_107_429 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_107_441 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_107_447 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_107_449 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_107_461 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_107_473 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_107_485 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_107_497 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_107_503 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_8 FILLER_107_505 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_4 FILLER_107_51 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_107_513 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_107_55 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_107_57 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_107_69 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_107_81 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_107_93 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_108_109 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_108_121 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_108_133 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_108_139 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_108_141 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_108_15 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_108_153 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_108_165 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_108_177 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_108_189 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_108_195 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_108_197 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_108_209 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_108_221 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_108_233 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_108_245 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_108_251 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_108_253 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_108_265 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_108_27 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_108_277 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_108_289 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_108_29 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_108_3 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_108_301 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_108_307 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_108_309 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_108_321 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_108_333 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_108_345 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_108_357 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_108_363 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_108_365 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_108_377 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_108_389 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_108_401 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_108_41 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_108_413 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_108_419 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_108_421 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_108_433 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_108_445 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_108_457 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_108_469 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_108_475 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_108_477 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_108_489 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_108_501 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_108_513 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_108_53 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_108_65 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_108_77 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_108_83 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_108_85 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_108_97 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_109_105 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_109_111 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_109_113 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_109_125 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_109_137 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_109_149 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_109_15 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_109_161 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_109_167 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_109_169 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_109_181 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_109_193 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_109_205 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_109_217 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_109_223 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_109_225 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_109_237 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_109_249 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_109_261 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_109_27 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_109_273 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_109_279 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_109_281 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_109_293 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_109_3 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_109_305 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_109_317 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_109_329 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_109_335 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_109_337 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_109_349 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_109_361 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_109_373 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_109_385 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_109_39 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_109_391 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_109_393 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_109_405 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_109_417 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_109_429 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_109_441 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_109_447 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_109_449 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_109_461 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_109_473 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_109_485 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_109_497 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_109_503 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_8 FILLER_109_505 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_4 FILLER_109_51 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_109_513 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_109_55 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_109_57 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_109_69 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_109_81 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_109_93 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_10_109 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_10_121 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_10_133 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_10_139 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_10_141 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_10_15 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_10_153 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_10_165 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_10_177 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_10_189 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_10_195 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_10_197 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_10_209 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_10_221 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_10_233 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_10_245 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_10_251 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_10_253 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_10_265 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_10_27 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_10_277 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_10_289 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_10_29 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_10_3 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_10_301 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_10_307 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_10_309 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_10_321 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_10_333 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_10_345 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_10_357 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_10_363 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_10_365 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_10_377 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_10_389 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_10_401 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_10_41 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_10_413 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_10_419 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_10_421 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_10_433 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_10_445 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_10_457 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_10_469 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_10_475 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_10_477 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_10_489 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_10_501 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_10_513 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_10_53 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_10_65 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_10_77 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_10_83 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_10_85 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_10_97 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_110_109 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_110_121 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_110_133 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_110_139 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_110_141 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_110_15 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_110_153 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_110_165 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_110_177 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_110_189 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_110_195 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_110_197 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_110_209 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_110_221 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_110_233 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_110_245 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_110_251 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_110_253 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_110_265 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_110_27 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_110_277 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_110_289 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_110_29 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_110_3 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_110_301 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_110_307 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_110_309 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_110_321 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_110_333 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_110_345 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_110_357 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_110_363 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_110_365 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_110_377 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_110_389 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_110_401 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_110_41 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_110_413 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_110_419 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_110_421 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_110_433 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_110_445 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_110_457 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_110_469 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_110_475 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_110_477 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_110_489 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_110_501 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_110_513 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_110_53 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_110_65 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_110_77 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_110_83 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_110_85 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_110_97 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_111_105 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_111_111 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_111_113 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_111_125 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_111_137 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_111_149 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_111_15 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_111_161 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_111_167 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_111_169 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_111_181 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_111_193 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_111_205 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_111_217 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_111_223 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_111_225 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_111_237 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_111_249 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_111_261 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_111_27 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_111_273 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_111_279 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_111_281 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_111_293 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_111_3 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_111_305 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_111_317 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_111_329 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_111_335 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_111_337 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_111_349 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_111_361 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_111_373 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_111_385 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_111_39 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_111_391 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_111_393 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_111_405 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_111_417 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_111_429 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_111_441 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_111_447 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_111_449 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_111_461 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_111_473 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_111_485 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_111_497 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_111_503 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_8 FILLER_111_505 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_4 FILLER_111_51 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_111_513 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_111_55 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_111_57 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_111_69 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_111_81 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_111_93 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_112_109 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_112_121 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_112_133 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_112_139 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_112_141 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_112_15 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_112_153 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_112_165 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_112_177 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_112_189 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_112_195 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_112_197 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_112_209 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_112_221 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_112_233 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_112_245 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_112_251 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_112_253 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_112_265 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_112_27 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_112_277 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_112_289 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_112_29 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_112_3 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_112_301 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_112_307 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_112_309 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_112_321 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_112_333 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_112_345 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_112_357 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_112_363 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_112_365 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_112_377 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_112_389 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_112_401 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_112_41 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_112_413 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_112_419 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_112_421 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_112_433 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_112_445 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_112_457 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_112_469 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_112_475 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_112_477 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_112_489 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_112_501 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_112_513 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_112_53 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_112_65 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_112_77 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_112_83 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_112_85 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_112_97 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_113_105 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_113_111 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_113_113 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_113_125 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_113_137 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_113_149 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_113_15 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_113_161 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_113_167 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_113_169 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_113_181 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_113_193 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_113_205 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_113_217 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_113_223 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_113_225 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_113_237 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_113_249 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_113_261 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_113_27 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_113_273 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_113_279 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_113_281 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_113_293 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_113_3 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_113_305 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_113_317 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_113_329 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_113_335 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_113_337 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_113_349 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_113_361 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_113_373 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_113_385 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_113_39 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_113_391 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_113_393 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_113_405 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_113_417 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_113_429 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_113_441 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_113_447 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_113_449 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_113_461 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_113_473 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_113_485 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_113_497 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_113_503 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_8 FILLER_113_505 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_4 FILLER_113_51 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_113_513 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_113_55 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_113_57 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_113_69 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_113_81 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_113_93 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_114_109 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_114_121 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_114_133 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_114_139 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_114_141 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_114_15 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_114_153 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_114_165 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_114_177 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_114_189 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_114_195 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_114_197 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_114_209 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_114_221 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_114_233 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_114_245 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_114_251 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_114_253 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_114_265 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_114_27 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_114_277 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_114_289 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_114_29 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_114_3 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_114_301 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_114_307 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_114_309 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_114_321 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_114_333 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_114_345 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_114_357 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_114_363 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_114_365 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_114_377 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_114_389 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_114_401 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_114_41 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_114_413 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_114_419 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_114_421 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_114_433 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_114_445 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_114_457 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_114_469 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_114_475 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_114_477 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_114_489 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_114_501 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_114_513 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_114_53 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_114_65 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_114_77 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_114_83 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_114_85 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_114_97 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_115_105 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_115_111 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_115_113 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_115_125 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_115_137 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_115_149 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_115_15 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_115_161 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_115_167 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_115_169 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_115_181 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_115_193 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_115_205 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_115_217 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_115_223 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_115_225 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_115_237 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_115_249 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_115_261 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_115_27 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_115_273 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_115_279 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_115_281 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_115_293 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_115_3 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_115_305 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_115_317 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_115_329 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_115_335 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_115_337 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_115_349 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_115_361 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_115_373 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_115_385 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_115_39 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_115_391 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_115_393 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_115_405 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_115_417 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_115_429 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_115_441 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_115_447 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_115_449 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_115_461 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_115_473 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_115_485 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_115_497 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_115_503 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_8 FILLER_115_505 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_4 FILLER_115_51 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_115_513 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_115_55 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_115_57 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_115_69 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_115_81 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_115_93 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_116_109 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_116_121 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_116_133 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_116_139 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_116_141 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_116_15 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_116_153 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_116_165 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_116_177 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_116_189 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_116_195 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_116_197 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_116_209 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_116_221 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_116_233 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_116_245 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_116_251 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_116_253 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_116_265 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_116_27 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_116_277 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_116_289 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_116_29 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_116_3 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_116_301 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_116_307 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_116_309 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_116_321 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_116_333 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_116_345 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_116_357 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_116_363 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_116_365 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_116_377 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_116_389 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_116_401 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_116_41 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_116_413 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_116_419 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_116_421 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_116_433 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_116_445 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_116_457 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_116_469 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_116_475 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_116_477 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_116_489 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_116_501 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_116_513 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_116_53 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_116_65 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_116_77 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_116_83 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_116_85 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_116_97 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_117_105 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_117_111 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_117_113 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_117_125 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_117_137 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_117_149 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_117_15 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_117_161 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_117_167 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_117_169 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_117_181 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_117_193 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_117_205 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_117_217 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_117_223 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_117_225 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_117_237 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_117_249 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_117_261 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_117_27 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_117_273 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_117_279 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_117_281 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_117_293 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_117_3 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_117_305 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_117_317 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_117_329 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_117_335 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_117_337 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_117_349 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_117_361 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_117_373 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_117_385 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_117_39 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_117_391 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_117_393 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_117_405 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_117_417 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_117_429 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_117_441 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_117_447 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_117_449 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_117_461 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_117_473 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_117_485 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_117_497 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_117_503 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_8 FILLER_117_505 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_4 FILLER_117_51 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_117_513 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_117_55 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_117_57 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_117_69 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_117_81 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_117_93 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_118_109 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_118_121 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_118_133 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_118_139 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_118_141 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_118_15 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_118_153 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_118_165 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_118_177 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_118_189 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_118_195 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_118_197 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_118_209 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_118_221 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_118_233 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_118_245 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_118_251 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_118_253 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_118_265 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_118_27 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_118_277 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_118_289 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_118_29 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_118_3 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_118_301 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_118_307 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_118_309 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_118_321 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_118_333 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_118_345 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_118_357 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_118_363 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_118_365 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_118_377 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_118_389 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_118_401 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_118_41 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_118_413 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_118_419 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_118_421 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_118_433 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_118_445 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_118_457 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_118_469 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_118_475 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_118_477 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_118_489 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_118_501 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_118_513 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_118_53 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_118_65 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_118_77 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_118_83 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_118_85 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_118_97 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_119_105 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_119_111 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_119_113 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_119_125 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_119_137 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_119_149 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_119_15 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_119_161 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_119_167 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_119_169 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_119_181 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_119_193 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_119_205 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_119_217 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_119_223 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_119_225 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_119_237 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_119_249 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_119_261 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_119_27 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_119_273 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_119_279 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_119_281 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_119_293 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_119_3 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_119_305 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_119_317 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_119_329 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_119_335 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_119_337 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_119_349 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_119_361 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_119_373 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_119_385 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_119_39 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_119_391 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_119_393 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_119_405 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_119_417 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_119_429 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_119_441 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_119_447 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_119_449 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_119_461 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_119_473 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_119_485 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_119_497 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_119_503 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_8 FILLER_119_505 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_4 FILLER_119_51 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_119_513 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_119_55 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_119_57 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_119_69 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_119_81 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_119_93 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_11_105 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_11_111 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_11_113 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_11_125 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_11_137 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_11_149 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_11_15 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_11_161 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_11_167 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_11_169 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_11_181 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_11_193 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_11_205 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_11_217 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_11_223 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_11_225 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_11_237 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_11_249 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_11_261 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_11_27 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_11_273 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_11_279 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_11_281 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_11_293 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_11_3 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_11_305 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_11_317 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_11_329 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_11_335 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_11_337 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_11_349 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_11_361 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_11_373 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_11_385 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_11_39 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_11_391 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_11_393 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_11_405 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_11_417 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_11_429 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_11_441 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_11_447 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_11_449 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_11_461 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_11_473 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_11_485 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_11_497 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_11_503 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_8 FILLER_11_505 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_4 FILLER_11_51 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_11_513 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_11_55 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_11_57 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_11_69 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_11_81 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_11_93 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_120_109 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_120_121 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_120_133 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_120_139 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_120_141 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_120_15 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_120_153 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_120_165 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_120_177 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_120_189 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_120_195 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_120_197 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_120_209 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_120_221 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_120_233 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_120_245 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_120_251 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_120_253 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_120_265 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_120_27 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_120_277 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_120_289 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_120_29 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_120_3 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_120_301 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_120_307 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_120_309 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_120_321 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_120_333 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_120_345 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_120_357 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_120_363 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_120_365 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_120_377 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_120_389 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_120_401 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_120_41 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_120_413 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_120_419 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_120_421 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_120_433 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_120_445 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_120_457 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_120_469 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_120_475 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_120_477 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_120_489 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_120_501 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_120_513 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_120_53 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_120_65 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_120_77 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_120_83 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_120_85 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_120_97 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_121_105 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_121_111 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_121_113 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_121_125 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_121_137 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_121_149 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_121_15 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_121_161 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_121_167 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_121_169 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_121_181 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_121_193 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_121_205 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_121_217 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_121_223 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_121_225 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_121_237 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_121_249 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_121_261 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_121_27 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_121_273 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_121_279 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_121_281 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_121_293 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_121_3 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_121_305 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_121_317 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_121_329 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_121_335 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_121_337 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_121_349 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_121_361 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_121_373 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_121_385 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_121_39 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_121_391 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_121_393 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_121_405 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_121_417 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_121_429 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_121_441 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_121_447 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_121_449 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_121_461 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_121_473 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_121_485 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_121_497 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_121_503 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_8 FILLER_121_505 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_4 FILLER_121_51 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_121_513 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_121_55 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_121_57 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_121_69 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_121_81 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_121_93 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_122_109 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_122_121 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_122_133 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_122_139 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_122_141 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_122_15 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_122_153 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_122_165 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_122_177 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_122_189 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_122_195 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_122_197 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_122_209 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_122_221 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_122_233 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_122_245 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_122_251 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_122_253 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_122_265 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_122_27 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_122_277 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_122_289 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_122_29 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_122_3 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_122_301 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_122_307 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_122_309 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_122_321 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_122_333 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_122_345 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_122_357 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_122_363 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_122_365 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_122_377 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_122_389 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_122_401 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_122_41 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_122_413 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_122_419 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_122_421 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_122_433 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_122_445 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_122_457 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_122_469 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_122_475 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_122_477 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_122_489 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_122_501 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_122_513 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_122_53 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_122_65 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_122_77 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_122_83 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_122_85 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_122_97 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_123_105 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_123_111 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_123_113 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_123_125 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_123_137 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_123_149 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_123_15 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_123_161 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_123_167 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_123_169 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_123_181 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_123_193 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_123_205 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_123_217 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_123_223 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_123_225 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_123_237 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_123_249 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_123_261 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_123_27 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_123_273 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_123_279 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_123_281 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_123_293 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_123_3 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_123_305 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_123_317 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_123_329 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_123_335 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_123_337 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_123_349 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_123_361 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_123_373 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_123_385 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_123_39 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_123_391 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_123_393 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_123_405 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_123_417 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_123_429 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_123_441 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_123_447 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_123_449 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_123_461 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_123_473 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_123_485 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_123_497 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_123_503 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_8 FILLER_123_505 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_4 FILLER_123_51 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_123_513 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_123_55 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_123_57 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_123_69 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_123_81 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_123_93 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_124_109 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_124_121 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_124_133 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_124_139 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_124_141 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_124_15 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_124_153 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_124_165 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_124_177 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_124_189 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_124_195 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_124_197 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_124_209 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_124_221 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_124_233 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_124_245 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_124_251 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_124_253 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_124_265 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_124_27 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_124_277 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_124_289 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_124_29 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_124_3 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_124_301 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_124_307 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_124_309 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_124_321 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_124_333 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_124_345 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_124_357 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_124_363 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_124_365 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_124_377 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_124_389 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_124_401 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_124_41 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_124_413 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_124_419 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_124_421 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_124_433 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_124_445 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_124_457 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_124_469 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_124_475 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_124_477 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_124_489 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_124_501 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_124_513 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_124_53 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_124_65 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_124_77 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_124_83 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_124_85 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_124_97 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_125_105 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_125_111 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_125_113 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_125_125 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_125_137 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_125_149 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_125_15 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_125_161 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_125_167 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_125_169 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_125_181 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_125_193 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_125_205 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_125_217 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_125_223 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_125_225 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_125_237 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_125_249 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_125_261 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_125_27 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_125_273 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_125_279 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_125_281 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_125_293 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_125_3 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_125_305 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_125_317 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_125_329 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_125_335 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_125_337 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_125_349 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_125_361 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_125_373 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_125_385 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_125_39 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_125_391 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_125_393 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_125_405 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_125_417 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_125_429 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_125_441 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_125_447 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_125_449 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_125_461 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_125_473 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_125_485 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_125_497 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_125_503 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_8 FILLER_125_505 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_4 FILLER_125_51 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_125_513 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_125_55 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_125_57 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_125_69 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_125_81 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_125_93 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_126_109 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_126_121 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_126_133 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_126_139 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_126_141 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_126_15 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_126_153 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_126_165 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_126_177 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_126_189 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_126_195 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_126_197 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_126_209 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_126_221 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_126_233 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_126_245 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_126_251 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_126_253 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_126_265 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_126_27 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_126_277 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_126_289 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_126_29 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_126_3 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_126_301 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_126_307 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_126_309 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_126_321 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_126_333 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_126_345 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_126_357 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_126_363 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_126_365 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_126_377 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_126_389 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_126_401 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_126_41 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_126_413 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_126_419 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_126_421 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_126_433 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_126_445 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_126_457 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_126_469 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_126_475 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_126_477 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_126_489 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_126_501 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_126_513 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_126_53 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_126_65 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_126_77 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_126_83 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_126_85 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_126_97 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_127_105 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_127_111 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_127_113 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_127_125 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_127_137 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_127_149 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_127_15 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_127_161 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_127_167 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_127_169 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_127_181 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_127_193 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_127_205 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_127_217 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_127_223 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_127_225 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_127_237 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_127_249 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_127_261 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_127_27 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_127_273 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_127_279 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_127_281 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_127_293 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_127_3 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_127_305 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_127_317 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_127_329 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_127_335 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_127_337 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_127_349 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_127_361 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_127_373 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_127_385 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_127_39 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_127_391 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_127_393 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_127_405 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_127_417 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_127_429 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_127_441 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_127_447 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_127_449 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_127_461 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_127_473 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_127_485 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_127_497 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_127_503 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_8 FILLER_127_505 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_4 FILLER_127_51 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_127_513 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_127_55 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_127_57 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_127_69 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_127_81 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_127_93 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_128_109 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_128_121 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_128_133 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_128_139 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_128_141 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_128_15 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_128_153 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_128_165 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_128_177 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_128_189 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_128_195 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_128_197 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_128_209 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_128_221 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_128_233 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_128_245 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_128_251 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_128_253 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_128_265 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_128_27 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_128_277 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_128_289 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_128_29 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_128_3 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_128_301 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_128_307 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_128_309 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_128_321 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_128_333 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_128_345 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_128_357 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_128_363 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_128_365 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_128_377 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_128_389 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_128_401 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_128_41 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_128_413 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_128_419 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_128_421 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_128_433 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_128_445 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_128_457 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_128_469 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_128_475 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_128_477 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_128_489 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_128_501 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_128_513 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_128_53 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_128_65 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_128_77 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_128_83 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_128_85 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_128_97 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_129_105 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_129_111 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_129_113 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_129_125 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_129_137 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_129_149 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_129_15 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_129_161 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_129_167 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_129_169 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_129_181 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_129_193 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_129_205 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_129_217 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_129_223 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_129_225 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_129_237 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_129_249 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_129_261 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_129_27 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_129_273 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_129_279 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_129_281 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_129_293 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_129_3 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_129_305 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_129_317 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_129_329 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_129_335 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_129_337 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_129_349 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_129_361 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_129_373 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_129_385 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_129_39 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_129_391 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_129_393 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_129_405 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_129_417 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_129_429 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_129_441 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_129_447 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_129_449 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_129_461 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_129_473 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_129_485 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_129_497 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_129_503 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_8 FILLER_129_505 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_4 FILLER_129_51 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_129_513 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_129_55 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_129_57 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_129_69 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_129_81 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_129_93 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_12_109 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_12_121 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_12_133 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_12_139 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_12_141 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_12_15 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_12_153 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_12_165 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_12_177 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_12_189 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_12_195 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_12_197 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_12_209 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_12_221 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_12_233 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_12_245 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_12_251 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_12_253 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_12_265 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_12_27 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_12_277 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_12_289 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_12_29 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_12_3 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_12_301 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_12_307 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_12_309 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_12_321 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_12_333 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_12_345 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_12_357 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_12_363 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_12_365 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_12_377 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_12_389 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_12_401 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_12_41 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_12_413 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_12_419 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_12_421 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_12_433 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_12_445 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_12_457 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_12_469 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_12_475 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_12_477 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_12_489 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_12_501 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_12_513 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_12_53 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_12_65 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_12_77 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_12_83 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_12_85 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_12_97 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_130_109 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_130_121 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_130_133 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_130_139 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_130_141 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_130_15 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_130_153 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_130_165 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_130_177 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_130_189 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_130_195 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_130_197 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_130_209 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_130_221 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_130_233 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_130_245 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_130_251 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_130_253 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_130_265 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_130_27 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_130_277 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_130_289 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_130_29 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_130_3 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_130_301 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_130_307 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_130_309 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_130_321 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_130_333 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_130_345 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_130_357 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_130_363 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_130_365 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_130_377 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_130_389 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_130_401 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_130_41 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_130_413 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_130_419 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_130_421 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_130_433 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_130_445 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_130_457 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_130_469 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_130_475 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_130_477 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_130_489 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_130_501 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_130_513 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_130_53 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_130_65 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_130_77 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_130_83 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_130_85 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_130_97 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_131_105 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_131_111 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_131_113 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_131_125 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_131_137 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_131_149 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_131_15 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_131_161 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_131_167 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_131_169 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_131_181 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_131_193 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_131_205 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_131_217 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_131_223 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_131_225 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_131_237 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_131_249 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_131_261 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_131_27 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_131_273 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_131_279 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_131_281 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_131_293 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_131_3 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_131_305 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_131_317 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_131_329 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_131_335 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_131_337 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_131_349 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_131_361 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_131_373 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_131_385 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_131_39 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_131_391 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_131_393 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_131_405 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_131_417 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_131_429 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_131_441 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_131_447 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_131_449 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_131_461 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_131_473 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_131_485 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_131_497 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_131_503 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_8 FILLER_131_505 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_4 FILLER_131_51 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_131_513 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_131_55 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_131_57 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_131_69 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_131_81 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_131_93 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_132_109 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_132_121 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_132_133 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_132_139 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_132_141 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_132_15 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_132_153 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_132_165 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_132_177 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_132_189 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_132_195 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_132_197 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_132_209 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_132_221 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_132_233 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_132_245 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_132_251 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_132_253 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_132_265 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_132_27 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_132_277 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_132_289 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_132_29 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_132_3 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_132_301 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_132_307 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_132_309 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_132_321 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_132_333 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_132_345 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_132_357 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_132_363 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_132_365 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_132_377 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_132_389 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_132_401 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_132_41 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_132_413 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_132_419 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_132_421 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_132_433 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_132_445 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_132_457 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_132_469 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_132_475 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_132_477 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_132_489 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_132_501 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_132_513 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_132_53 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_132_65 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_132_77 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_132_83 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_132_85 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_132_97 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_133_105 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_133_111 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_133_113 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_133_125 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_133_137 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_133_149 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_133_15 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_133_161 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_133_167 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_133_169 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_133_181 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_133_193 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_133_205 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_133_217 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_133_223 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_133_225 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_133_237 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_133_249 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_133_261 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_133_27 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_133_273 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_133_279 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_133_281 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_133_293 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_133_3 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_133_305 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_133_317 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_133_329 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_133_335 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_133_337 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_133_349 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_133_361 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_133_373 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_133_385 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_133_39 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_133_391 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_133_393 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_133_405 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_133_417 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_133_429 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_133_441 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_133_447 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_133_449 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_133_461 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_133_473 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_133_485 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_133_497 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_133_503 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_8 FILLER_133_505 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_4 FILLER_133_51 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_133_513 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_133_55 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_133_57 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_133_69 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_133_81 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_133_93 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_134_109 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_134_121 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_134_133 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_134_139 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_134_141 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_134_15 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_134_153 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_134_165 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_134_177 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_134_189 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_134_195 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_134_197 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_134_209 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_134_221 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_134_233 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_134_245 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_134_251 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_134_253 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_134_265 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_134_27 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_134_277 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_134_289 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_134_29 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_134_3 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_134_301 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_134_307 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_134_309 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_134_321 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_134_333 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_134_345 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_134_357 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_134_363 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_134_365 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_134_377 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_134_389 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_134_401 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_134_41 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_134_413 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_134_419 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_134_421 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_134_433 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_134_445 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_134_457 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_134_469 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_134_475 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_134_477 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_134_489 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_134_501 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_134_513 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_134_53 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_134_65 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_134_77 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_134_83 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_134_85 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_134_97 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_135_105 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_135_111 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_135_113 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_135_125 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_135_137 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_135_149 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_135_15 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_135_161 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_135_167 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_135_169 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_135_181 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_135_193 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_135_205 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_135_217 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_135_223 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_135_225 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_135_237 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_135_249 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_135_261 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_135_27 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_135_273 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_135_279 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_135_281 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_135_293 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_135_3 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_135_305 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_135_317 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_135_329 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_135_335 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_135_337 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_135_349 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_135_361 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_135_373 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_135_385 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_135_39 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_135_391 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_135_393 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_135_405 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_135_417 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_135_429 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_135_441 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_135_447 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_135_449 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_135_461 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_135_473 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_135_485 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_135_497 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_135_503 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_8 FILLER_135_505 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_4 FILLER_135_51 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_135_513 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_135_55 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_135_57 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_135_69 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_135_81 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_135_93 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_136_109 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_136_121 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_136_133 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_136_139 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_136_141 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_136_15 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_136_153 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_136_165 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_136_177 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_136_189 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_136_195 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_136_197 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_136_209 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_136_221 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_136_233 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_136_245 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_136_251 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_136_253 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_136_265 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_136_27 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_136_277 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_136_289 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_136_29 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_136_3 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_136_301 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_136_307 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_136_309 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_136_321 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_136_333 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_136_345 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_136_357 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_136_363 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_136_365 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_136_377 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_136_389 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_136_401 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_136_41 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_136_413 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_136_419 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_136_421 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_136_433 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_136_445 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_136_457 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_136_469 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_136_475 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_136_477 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_136_489 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_136_501 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_136_513 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_136_53 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_136_65 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_136_77 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_136_83 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_136_85 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_136_97 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_137_105 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_137_111 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_137_113 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_137_125 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_137_137 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_137_149 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_137_15 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_137_161 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_137_167 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_137_169 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_137_181 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_137_193 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_137_205 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_137_217 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_137_223 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_137_225 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_137_237 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_137_249 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_137_261 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_137_27 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_137_273 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_137_279 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_137_281 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_137_293 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_137_3 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_137_305 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_137_317 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_137_329 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_137_335 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_137_337 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_137_349 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_137_361 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_137_373 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_137_385 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_137_39 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_137_391 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_137_393 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_137_405 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_137_417 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_137_429 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_137_441 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_137_447 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_137_449 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_137_461 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_137_473 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_137_485 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_137_497 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_137_503 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_8 FILLER_137_505 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_4 FILLER_137_51 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_137_513 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_137_55 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_137_57 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_137_69 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_137_81 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_137_93 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_138_109 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_138_121 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_138_133 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_138_139 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_138_141 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_138_15 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_138_153 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_138_165 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_138_177 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_138_189 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_138_195 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_138_197 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_138_209 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_138_221 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_138_233 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_138_245 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_138_251 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_138_253 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_138_265 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_138_27 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_138_277 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_138_289 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_138_29 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_138_3 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_138_301 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_138_307 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_138_309 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_138_321 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_138_333 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_138_345 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_138_357 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_138_363 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_138_365 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_138_377 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_138_389 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_138_401 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_138_41 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_138_413 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_138_419 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_138_421 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_138_433 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_138_445 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_138_457 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_138_469 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_138_475 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_138_477 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_138_489 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_138_501 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_138_513 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_138_53 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_138_65 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_138_77 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_138_83 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_138_85 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_138_97 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_139_105 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_139_111 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_139_113 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_139_125 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_139_137 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_139_149 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_139_15 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_139_161 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_139_167 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_139_169 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_139_181 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_139_193 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_139_205 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_139_217 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_139_223 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_139_225 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_139_237 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_139_249 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_139_261 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_139_27 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_139_273 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_139_279 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_139_281 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_139_293 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_139_3 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_139_305 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_139_317 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_139_329 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_139_335 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_139_337 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_139_349 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_139_361 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_139_373 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_139_385 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_139_39 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_139_391 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_139_393 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_139_405 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_139_417 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_139_429 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_139_441 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_139_447 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_139_449 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_139_461 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_139_473 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_139_485 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_139_497 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_139_503 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_8 FILLER_139_505 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_4 FILLER_139_51 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_139_513 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_139_55 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_139_57 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_139_69 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_139_81 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_139_93 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_13_105 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_13_111 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_13_113 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_13_125 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_13_137 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_13_149 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_13_15 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_13_161 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_13_167 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_13_169 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_13_181 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_13_193 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_13_205 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_13_217 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_13_223 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_13_225 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_13_237 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_13_249 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_13_261 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_13_27 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_13_273 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_13_279 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_13_281 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_13_293 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_13_3 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_13_305 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_13_317 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_13_329 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_13_335 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_13_337 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_13_349 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_13_361 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_13_373 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_13_385 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_13_39 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_13_391 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_13_393 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_13_405 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_13_417 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_13_429 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_13_441 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_13_447 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_13_449 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_13_461 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_13_473 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_13_485 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_13_497 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_13_503 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_8 FILLER_13_505 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_4 FILLER_13_51 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_13_513 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_13_55 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_13_57 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_13_69 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_13_81 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_13_93 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_140_109 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_140_121 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_140_133 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_140_139 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_140_141 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_140_15 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_140_153 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_140_165 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_140_177 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_140_189 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_140_195 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_140_197 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_140_209 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_140_221 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_140_233 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_140_245 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_140_251 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_140_253 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_140_265 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_140_27 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_140_277 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_140_289 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_140_29 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_140_3 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_140_301 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_140_307 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_140_309 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_140_321 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_140_333 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_140_345 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_140_357 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_140_363 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_140_365 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_140_377 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_140_389 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_140_401 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_140_41 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_140_413 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_140_419 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_140_421 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_140_433 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_140_445 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_140_457 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_140_469 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_140_475 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_140_477 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_140_489 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_140_501 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_140_513 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_140_53 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_140_65 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_140_77 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_140_83 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_140_85 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_140_97 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_141_105 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_141_111 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_141_113 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_141_125 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_141_137 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_141_149 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_141_15 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_141_161 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_141_167 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_141_169 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_141_181 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_141_193 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_141_205 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_141_217 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_141_223 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_141_225 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_141_237 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_141_249 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_141_261 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_141_27 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_141_273 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_141_279 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_141_281 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_141_293 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_141_3 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_141_305 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_141_317 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_141_329 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_141_335 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_141_337 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_141_349 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_141_361 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_141_373 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_141_385 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_141_39 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_141_391 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_141_393 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_141_405 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_141_417 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_141_429 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_141_441 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_141_447 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_141_449 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_141_461 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_141_473 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_141_485 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_141_497 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_141_503 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_8 FILLER_141_505 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_4 FILLER_141_51 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_141_513 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_141_55 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_141_57 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_141_69 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_141_81 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_141_93 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_142_109 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_142_121 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_142_133 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_142_139 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_142_141 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_142_15 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_142_153 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_142_165 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_142_177 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_142_189 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_142_195 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_142_197 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_142_209 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_142_221 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_142_233 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_142_245 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_142_251 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_142_253 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_142_265 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_142_27 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_142_277 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_142_289 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_142_29 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_142_3 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_142_301 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_142_307 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_142_309 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_142_321 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_142_333 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_142_345 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_142_357 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_142_363 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_142_365 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_142_377 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_142_389 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_142_401 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_142_41 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_142_413 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_142_419 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_142_421 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_142_433 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_142_445 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_142_457 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_142_469 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_142_475 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_142_477 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_142_489 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_142_501 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_142_513 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_142_53 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_142_65 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_142_77 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_142_83 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_142_85 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_142_97 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_143_105 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_143_111 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_143_113 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_143_125 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_143_137 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_143_149 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_143_15 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_143_161 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_143_167 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_143_169 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_143_181 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_143_193 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_143_205 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_143_217 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_143_223 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_143_225 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_143_237 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_143_249 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_143_261 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_143_27 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_143_273 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_143_279 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_143_281 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_143_293 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_143_3 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_143_305 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_143_317 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_143_329 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_143_335 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_143_337 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_143_349 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_143_361 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_143_373 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_143_385 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_143_39 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_143_391 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_143_393 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_143_405 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_143_417 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_143_429 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_143_441 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_143_447 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_143_449 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_143_461 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_143_473 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_143_485 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_143_497 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_143_503 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_8 FILLER_143_505 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_4 FILLER_143_51 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_143_513 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_143_55 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_143_57 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_143_69 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_143_81 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_143_93 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_144_109 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_144_121 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_144_133 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_144_139 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_144_141 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_144_15 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_144_153 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_144_165 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_144_177 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_144_189 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_144_195 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_144_197 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_144_209 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_144_221 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_144_233 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_144_245 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_144_251 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_144_253 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_144_265 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_144_27 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_144_277 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_144_289 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_144_29 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_144_3 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_144_301 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_144_307 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_144_309 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_144_321 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_144_333 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_144_345 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_144_357 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_144_363 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_144_365 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_144_377 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_144_389 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_144_401 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_144_41 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_144_413 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_144_419 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_144_421 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_144_433 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_144_445 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_144_457 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_144_469 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_144_475 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_144_477 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_144_489 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_144_501 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_144_513 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_144_53 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_144_65 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_144_77 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_144_83 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_144_85 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_144_97 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_145_105 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_145_111 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_145_113 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_145_125 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_145_137 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_145_149 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_145_15 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_145_161 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_145_167 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_145_169 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_145_181 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_145_193 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_145_205 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_145_217 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_145_223 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_145_225 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_145_237 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_145_249 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_145_261 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_145_27 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_145_273 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_145_279 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_145_281 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_145_293 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_145_3 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_145_305 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_145_317 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_145_329 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_145_335 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_145_337 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_145_349 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_145_361 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_145_373 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_145_385 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_145_39 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_145_391 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_145_393 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_145_405 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_145_417 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_145_429 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_145_441 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_145_447 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_145_449 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_145_461 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_145_473 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_145_485 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_145_497 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_145_503 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_8 FILLER_145_505 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_4 FILLER_145_51 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_145_513 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_145_55 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_145_57 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_145_69 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_145_81 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_145_93 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_146_109 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_146_121 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_146_133 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_146_139 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_146_141 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_146_15 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_146_153 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_146_165 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_146_177 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_146_189 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_146_195 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_146_197 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_146_209 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_146_221 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_146_233 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_146_245 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_146_251 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_146_253 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_146_265 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_146_27 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_146_277 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_146_289 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_146_29 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_146_3 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_146_301 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_146_307 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_146_309 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_146_321 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_146_333 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_146_345 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_146_357 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_146_363 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_146_365 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_146_377 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_146_389 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_146_401 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_146_41 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_146_413 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_146_419 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_146_421 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_146_433 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_146_445 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_146_457 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_146_469 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_146_475 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_146_477 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_146_489 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_146_501 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_146_513 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_146_53 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_146_65 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_146_77 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_146_83 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_146_85 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_146_97 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_147_105 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_147_111 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_147_113 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_147_125 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_147_137 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_147_149 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_147_15 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_147_161 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_147_167 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_147_169 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_147_181 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_147_193 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_147_205 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_147_217 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_147_223 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_147_225 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_147_237 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_147_249 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_147_261 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_147_27 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_147_273 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_147_279 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_147_281 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_147_293 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_147_3 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_147_305 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_147_317 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_147_329 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_147_335 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_147_337 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_147_349 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_147_361 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_147_373 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_147_385 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_147_39 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_147_391 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_147_393 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_147_405 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_147_417 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_147_429 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_147_441 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_147_447 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_147_449 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_147_461 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_147_473 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_147_485 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_147_497 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_147_503 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_8 FILLER_147_505 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_4 FILLER_147_51 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_147_513 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_147_55 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_147_57 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_147_69 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_147_81 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_147_93 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_148_109 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_148_121 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_148_133 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_148_139 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_148_141 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_148_15 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_148_153 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_148_165 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_148_177 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_148_189 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_148_195 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_148_197 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_148_209 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_148_221 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_148_233 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_148_245 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_148_251 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_148_253 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_148_265 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_148_27 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_148_277 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_148_289 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_148_29 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_148_3 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_148_301 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_148_307 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_148_309 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_148_321 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_148_333 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_148_345 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_148_357 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_148_363 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_148_365 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_148_377 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_148_389 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_148_401 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_148_41 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_148_413 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_148_419 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_148_421 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_148_433 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_148_445 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_148_457 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_148_469 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_148_475 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_148_477 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_148_489 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_148_501 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_148_513 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_148_53 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_148_65 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_148_77 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_148_83 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_148_85 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_148_97 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_149_105 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_149_111 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_149_113 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_149_125 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_149_137 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_149_149 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_149_15 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_149_161 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_149_167 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_149_169 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_149_181 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_149_193 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_149_205 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_149_217 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_149_223 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_149_225 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_149_237 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_149_249 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_149_261 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_149_27 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_149_273 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_149_279 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_149_281 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_149_293 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_149_3 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_149_305 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_149_317 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_149_329 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_149_335 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_149_337 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_149_349 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_149_361 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_149_373 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_149_385 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_149_39 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_149_391 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_149_393 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_149_405 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_149_417 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_149_429 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_149_441 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_149_447 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_149_449 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_149_461 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_149_473 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_149_485 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_149_497 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_149_503 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_8 FILLER_149_505 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_4 FILLER_149_51 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_149_513 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_149_55 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_149_57 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_149_69 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_149_81 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_149_93 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_14_109 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_14_121 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_14_133 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_14_139 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_14_141 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_14_15 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_14_153 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_14_165 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_14_177 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_14_189 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_14_195 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_14_197 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_14_209 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_14_221 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_14_233 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_14_245 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_14_251 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_14_253 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_14_265 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_14_27 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_14_277 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_14_289 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_14_29 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_14_3 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_14_301 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_14_307 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_14_309 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_14_321 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_14_333 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_14_345 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_14_357 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_14_363 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_14_365 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_14_377 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_14_389 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_14_401 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_14_41 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_14_413 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_14_419 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_14_421 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_14_433 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_14_445 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_14_457 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_14_469 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_14_475 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_14_477 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_14_489 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_14_501 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_14_513 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_14_53 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_14_65 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_14_77 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_14_83 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_14_85 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_14_97 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_150_109 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_150_121 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_150_133 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_150_139 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_150_141 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_150_15 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_150_153 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_150_165 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_150_177 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_150_189 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_150_195 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_150_197 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_150_209 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_150_221 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_150_233 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_150_245 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_150_251 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_150_253 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_150_265 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_150_27 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_150_277 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_150_289 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_150_29 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_150_3 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_150_301 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_150_307 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_150_309 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_150_321 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_150_333 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_150_345 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_150_357 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_150_363 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_150_365 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_150_377 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_150_389 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_150_401 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_150_41 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_150_413 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_150_419 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_150_421 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_150_433 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_150_445 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_150_457 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_150_469 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_150_475 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_150_477 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_150_489 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_150_501 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_150_513 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_150_53 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_150_65 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_150_77 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_150_83 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_150_85 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_150_97 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_151_105 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_151_111 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_151_113 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_151_125 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_151_137 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_151_149 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_151_15 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_151_161 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_151_167 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_151_169 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_151_181 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_151_193 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_151_205 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_151_217 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_151_223 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_151_225 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_151_237 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_151_249 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_151_261 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_151_27 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_151_273 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_151_279 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_151_281 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_151_293 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_151_3 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_151_305 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_151_317 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_151_329 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_151_335 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_151_337 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_151_349 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_151_361 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_151_373 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_151_385 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_151_39 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_151_391 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_151_393 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_151_405 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_151_417 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_151_429 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_151_441 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_151_447 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_151_449 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_151_461 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_151_473 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_151_485 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_151_497 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_151_503 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_8 FILLER_151_505 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_4 FILLER_151_51 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_151_513 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_151_55 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_151_57 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_151_69 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_151_81 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_151_93 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_152_109 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_152_121 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_152_133 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_152_139 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_152_141 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_152_15 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_152_153 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_152_165 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_152_177 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_152_189 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_152_195 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_152_197 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_152_209 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_152_221 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_152_233 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_152_245 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_152_251 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_152_253 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_152_265 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_152_27 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_152_277 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_152_289 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_152_29 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_152_3 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_152_301 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_152_307 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_152_309 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_152_321 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_152_333 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_152_345 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_152_357 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_152_363 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_152_365 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_152_377 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_152_389 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_152_401 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_152_41 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_152_413 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_152_419 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_152_421 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_152_433 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_152_445 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_152_457 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_152_469 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_152_475 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_152_477 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_152_489 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_152_501 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_152_513 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_152_53 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_152_65 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_152_77 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_152_83 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_152_85 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_152_97 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_153_105 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_153_111 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_153_113 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_153_125 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_153_137 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_153_149 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_153_15 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_153_161 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_153_167 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_153_169 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_153_181 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_153_193 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_153_205 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_153_217 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_153_223 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_153_225 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_153_237 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_153_249 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_153_261 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_153_27 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_153_273 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_153_279 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_153_281 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_153_293 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_153_3 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_153_305 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_153_317 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_153_329 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_153_335 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_153_337 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_153_349 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_153_361 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_153_373 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_153_385 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_153_39 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_153_391 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_153_393 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_153_405 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_153_417 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_153_429 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_153_441 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_153_447 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_153_449 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_153_461 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_153_473 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_153_485 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_153_497 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_153_503 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_8 FILLER_153_505 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_4 FILLER_153_51 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_153_513 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_153_55 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_153_57 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_153_69 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_153_81 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_153_93 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_154_109 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_154_121 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_154_133 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_154_139 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_154_141 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_154_15 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_154_153 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_154_165 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_154_177 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_154_189 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_154_195 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_154_197 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_154_209 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_154_221 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_154_233 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_154_245 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_154_251 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_154_253 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_154_265 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_154_27 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_154_277 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_154_289 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_154_29 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_154_3 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_154_301 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_154_307 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_154_309 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_154_321 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_154_333 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_154_345 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_154_357 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_154_363 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_154_365 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_154_377 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_154_389 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_154_401 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_154_41 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_154_413 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_154_419 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_154_421 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_154_433 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_154_445 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_154_457 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_154_469 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_154_475 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_154_477 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_154_489 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_154_501 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_154_513 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_154_53 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_154_65 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_154_77 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_154_83 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_154_85 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_154_97 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_155_105 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_155_111 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_155_113 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_155_125 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_155_137 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_155_149 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_155_15 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_155_161 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_155_167 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_155_169 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_155_181 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_155_193 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_155_205 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_155_217 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_155_223 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_155_225 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_155_237 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_155_249 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_155_261 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_155_27 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_155_273 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_155_279 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_155_281 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_155_293 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_155_3 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_155_305 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_155_317 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_155_329 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_155_335 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_155_337 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_155_349 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_155_361 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_155_373 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_155_385 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_155_39 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_155_391 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_155_393 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_155_405 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_155_417 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_155_429 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_155_441 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_155_447 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_155_449 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_155_461 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_155_473 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_155_485 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_155_497 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_155_503 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_8 FILLER_155_505 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_4 FILLER_155_51 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_155_513 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_155_55 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_155_57 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_155_69 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_155_81 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_155_93 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_156_109 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_156_121 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_156_133 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_156_139 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_156_141 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_156_15 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_156_153 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_156_165 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_156_177 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_156_189 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_156_195 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_156_197 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_156_209 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_156_221 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_156_233 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_156_245 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_156_251 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_156_253 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_156_265 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_156_27 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_156_277 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_156_289 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_156_29 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_156_3 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_156_301 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_156_307 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_156_309 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_156_321 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_156_333 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_156_345 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_156_357 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_156_363 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_156_365 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_156_377 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_156_389 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_156_401 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_156_41 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_156_413 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_156_419 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_156_421 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_156_433 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_156_445 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_156_457 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_156_469 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_156_475 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_156_477 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_156_489 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_156_501 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_156_513 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_156_53 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_156_65 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_156_77 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_156_83 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_156_85 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_156_97 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_157_105 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_157_111 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_157_113 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_157_125 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_157_137 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_157_149 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_157_15 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_157_161 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_157_167 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_157_169 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_157_181 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_157_193 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_157_205 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_157_217 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_157_223 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_157_225 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_157_237 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_157_249 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_157_261 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_157_27 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_157_273 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_157_279 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_157_281 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_157_293 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_157_3 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_157_305 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_157_317 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_157_329 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_157_335 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_157_337 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_157_349 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_157_361 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_157_373 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_157_385 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_157_39 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_157_391 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_157_393 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_157_405 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_157_417 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_157_429 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_157_441 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_157_447 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_157_449 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_157_461 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_157_473 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_157_485 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_157_497 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_157_503 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_8 FILLER_157_505 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_4 FILLER_157_51 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_157_513 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_157_55 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_157_57 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_157_69 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_157_81 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_157_93 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_158_109 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_158_121 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_158_133 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_158_139 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_158_141 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_158_15 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_158_153 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_158_165 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_158_177 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_158_189 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_158_195 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_158_197 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_158_209 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_158_221 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_158_233 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_158_245 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_158_251 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_158_253 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_158_265 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_158_27 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_158_277 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_158_289 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_158_29 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_158_3 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_158_301 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_158_307 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_158_309 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_158_321 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_158_333 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_158_345 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_158_357 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_158_363 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_158_365 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_158_377 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_158_389 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_158_401 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_158_41 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_158_413 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_158_419 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_158_421 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_158_433 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_158_445 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_158_457 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_158_469 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_158_475 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_158_477 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_158_489 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_158_501 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_158_513 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_158_53 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_158_65 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_158_77 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_158_83 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_158_85 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_158_97 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_159_105 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_159_111 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_159_113 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_159_125 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_159_137 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_159_149 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_159_15 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_159_161 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_159_167 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_159_169 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_159_181 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_159_193 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_159_205 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_159_217 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_159_223 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_159_225 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_159_237 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_159_249 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_159_261 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_159_27 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_159_273 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_159_279 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_159_281 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_159_293 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_159_3 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_159_305 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_159_317 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_159_329 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_159_335 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_159_337 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_159_349 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_159_361 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_159_373 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_159_385 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_159_39 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_159_391 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_159_393 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_159_405 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_159_417 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_159_429 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_159_441 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_159_447 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_159_449 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_159_461 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_159_473 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_159_485 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_159_497 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_159_503 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_8 FILLER_159_505 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_4 FILLER_159_51 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_159_513 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_159_55 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_159_57 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_159_69 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_159_81 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_159_93 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_15_105 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_15_111 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_15_113 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_15_125 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_15_137 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_15_149 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_15_15 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_15_161 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_15_167 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_15_169 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_15_181 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_15_193 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_15_205 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_15_217 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_15_223 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_15_225 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_15_237 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_15_249 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_15_261 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_15_27 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_15_273 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_15_279 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_15_281 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_15_293 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_15_3 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_15_305 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_15_317 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_15_329 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_15_335 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_15_337 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_15_349 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_15_361 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_15_373 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_15_385 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_15_39 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_15_391 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_15_393 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_15_405 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_15_417 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_15_429 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_15_441 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_15_447 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_15_449 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_15_461 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_15_473 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_15_485 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_15_497 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_15_503 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_8 FILLER_15_505 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_4 FILLER_15_51 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_15_513 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_15_55 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_15_57 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_15_69 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_15_81 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_15_93 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_160_109 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_160_121 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_160_133 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_160_139 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_160_141 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_160_15 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_160_153 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_160_165 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_160_177 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_160_189 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_160_195 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_160_197 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_160_209 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_160_221 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_160_233 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_160_245 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_160_251 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_160_253 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_160_265 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_160_27 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_160_277 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_160_289 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_160_29 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_160_3 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_160_301 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_160_307 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_160_309 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_160_321 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_160_333 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_160_345 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_160_357 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_160_363 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_160_365 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_160_377 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_160_389 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_160_401 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_160_41 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_160_413 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_160_419 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_160_421 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_160_433 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_160_445 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_160_457 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_160_469 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_160_475 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_160_477 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_160_489 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_160_501 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_160_513 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_160_53 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_160_65 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_160_77 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_160_83 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_160_85 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_160_97 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_161_105 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_161_111 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_161_113 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_161_125 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_161_137 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_161_149 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_161_15 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_161_161 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_161_167 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_161_169 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_161_181 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_161_193 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_161_205 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_161_217 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_161_223 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_161_225 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_161_237 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_161_249 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_161_261 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_161_27 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_161_273 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_161_279 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_161_281 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_161_293 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_161_3 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_161_305 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_161_317 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_161_329 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_161_335 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_161_337 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_161_349 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_161_361 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_161_373 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_161_385 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_161_39 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_161_391 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_161_393 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_161_405 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_161_417 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_161_429 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_161_441 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_161_447 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_161_449 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_161_461 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_161_473 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_161_485 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_161_497 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_161_503 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_8 FILLER_161_505 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_4 FILLER_161_51 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_161_513 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_161_55 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_161_57 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_161_69 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_161_81 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_161_93 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_162_109 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_162_121 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_162_133 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_162_139 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_162_141 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_162_15 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_162_153 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_162_165 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_162_177 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_162_189 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_162_195 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_162_197 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_162_209 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_162_221 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_162_233 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_162_245 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_162_251 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_162_253 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_162_265 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_162_27 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_162_277 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_162_289 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_162_29 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_162_3 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_162_301 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_162_307 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_162_309 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_162_321 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_162_333 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_162_345 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_162_357 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_162_363 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_162_365 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_162_377 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_162_389 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_162_401 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_162_41 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_162_413 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_162_419 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_162_421 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_162_433 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_162_445 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_162_457 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_162_469 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_162_475 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_162_477 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_162_489 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_162_501 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_162_513 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_162_53 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_162_65 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_162_77 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_162_83 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_162_85 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_162_97 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_163_105 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_163_111 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_163_113 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_163_125 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_163_137 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_163_149 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_163_15 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_163_161 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_163_167 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_163_169 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_163_181 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_163_193 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_163_205 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_163_217 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_163_223 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_163_225 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_163_237 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_163_249 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_163_261 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_163_27 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_163_273 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_163_279 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_163_281 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_163_293 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_163_3 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_163_305 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_163_317 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_163_329 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_163_335 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_163_337 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_163_349 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_163_361 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_163_373 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_163_385 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_163_39 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_163_391 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_163_393 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_163_405 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_163_417 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_163_429 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_163_441 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_163_447 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_163_449 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_163_461 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_163_473 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_163_485 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_163_497 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_163_503 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_8 FILLER_163_505 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_4 FILLER_163_51 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_163_513 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_163_55 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_163_57 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_163_69 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_163_81 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_163_93 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_164_109 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_164_121 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_164_133 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_164_139 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_164_141 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_164_15 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_164_153 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_164_165 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_164_177 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_164_189 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_164_195 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_164_197 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_164_209 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_164_221 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_164_233 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_164_245 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_164_251 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_164_253 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_164_265 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_164_27 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_164_277 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_164_289 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_164_29 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_164_3 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_164_301 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_164_307 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_164_309 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_164_321 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_164_333 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_164_345 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_164_357 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_164_363 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_164_365 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_164_377 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_164_389 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_164_401 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_164_41 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_164_413 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_164_419 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_164_421 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_164_433 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_164_445 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_164_457 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_164_469 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_164_475 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_164_477 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_164_489 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_164_501 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_164_513 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_164_53 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_164_65 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_164_77 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_164_83 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_164_85 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_164_97 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_165_105 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_165_111 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_165_113 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_165_125 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_165_137 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_165_149 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_165_15 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_165_161 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_165_167 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_165_169 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_165_181 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_165_193 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_165_205 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_165_217 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_165_223 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_165_225 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_165_237 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_165_249 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_165_261 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_165_27 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_165_273 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_165_279 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_165_281 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_165_293 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_165_3 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_165_305 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_165_317 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_165_329 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_165_335 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_165_337 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_165_349 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_165_361 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_165_373 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_165_385 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_165_39 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_165_391 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_165_393 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_165_405 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_165_417 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_165_429 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_165_441 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_165_447 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_165_449 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_165_461 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_165_473 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_165_485 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_165_497 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_165_503 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_8 FILLER_165_505 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_4 FILLER_165_51 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_165_513 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_165_55 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_165_57 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_165_69 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_165_81 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_165_93 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_166_109 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_166_121 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_166_133 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_166_139 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_166_141 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_166_15 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_166_153 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_166_165 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_166_177 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_166_189 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_166_195 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_166_197 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_166_209 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_166_221 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_166_233 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_166_245 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_166_251 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_166_253 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_166_265 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_166_27 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_166_277 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_166_289 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_166_29 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_166_3 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_166_301 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_166_307 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_166_309 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_166_321 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_166_333 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_166_345 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_166_357 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_166_363 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_166_365 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_166_377 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_166_389 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_166_401 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_166_41 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_166_413 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_166_419 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_166_421 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_166_433 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_166_445 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_166_457 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_166_469 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_166_475 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_166_477 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_166_489 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_166_501 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_166_513 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_166_53 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_166_65 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_166_77 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_166_83 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_166_85 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_166_97 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_167_105 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_167_111 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_167_113 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_167_125 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_167_137 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_167_149 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_167_15 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_167_161 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_167_167 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_167_169 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_167_181 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_167_193 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_167_205 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_167_217 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_167_223 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_167_225 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_167_237 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_167_249 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_167_261 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_167_27 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_167_273 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_167_279 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_167_281 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_167_293 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_167_3 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_167_305 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_167_317 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_167_329 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_167_335 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_167_337 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_167_349 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_167_361 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_167_373 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_167_385 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_167_39 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_167_391 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_167_393 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_167_405 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_167_417 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_167_429 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_167_441 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_167_447 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_167_449 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_167_461 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_167_473 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_167_485 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_167_497 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_167_503 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_8 FILLER_167_505 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_4 FILLER_167_51 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_167_513 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_167_55 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_167_57 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_167_69 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_167_81 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_167_93 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_168_109 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_168_121 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_168_133 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_168_139 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_168_141 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_168_15 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_168_153 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_168_165 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_168_177 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_168_189 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_168_195 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_168_197 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_168_209 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_168_221 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_168_233 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_168_245 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_168_251 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_168_253 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_168_265 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_168_27 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_168_277 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_168_289 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_168_29 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_168_3 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_168_301 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_168_307 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_168_309 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_168_321 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_168_333 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_168_345 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_168_357 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_168_363 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_168_365 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_168_377 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_168_389 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_168_401 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_168_41 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_168_413 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_168_419 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_168_421 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_168_433 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_168_445 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_168_457 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_168_469 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_168_475 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_168_477 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_168_489 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_168_501 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_168_513 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_168_53 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_168_65 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_168_77 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_168_83 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_168_85 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_168_97 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_169_105 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_169_111 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_169_113 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_169_125 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_169_137 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_169_149 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_169_15 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_169_161 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_169_167 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_169_169 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_169_181 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_169_193 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_169_205 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_169_217 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_169_223 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_169_225 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_169_237 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_169_249 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_169_261 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_169_27 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_169_273 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_169_279 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_169_281 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_169_293 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_169_3 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_169_305 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_169_317 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_169_329 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_169_335 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_169_337 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_169_349 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_169_361 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_169_373 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_169_385 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_169_39 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_169_391 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_169_393 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_169_405 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_169_417 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_169_429 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_169_441 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_169_447 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_169_449 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_169_461 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_169_473 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_169_485 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_169_497 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_169_503 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_8 FILLER_169_505 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_4 FILLER_169_51 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_169_513 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_169_55 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_169_57 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_169_69 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_169_81 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_169_93 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_16_109 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_16_121 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_16_133 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_16_139 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_16_141 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_16_15 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_16_153 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_16_165 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_16_177 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_16_189 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_16_195 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_16_197 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_16_209 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_16_221 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_16_233 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_16_245 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_16_251 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_16_253 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_16_265 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_16_27 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_16_277 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_16_289 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_16_29 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_16_3 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_16_301 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_16_307 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_16_309 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_16_321 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_16_333 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_16_345 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_16_357 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_16_363 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_16_365 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_16_377 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_16_389 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_16_401 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_16_41 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_16_413 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_16_419 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_16_421 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_16_433 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_16_445 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_16_457 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_16_469 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_16_475 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_16_477 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_16_489 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_16_501 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_16_513 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_16_53 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_16_65 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_16_77 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_16_83 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_16_85 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_16_97 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_170_109 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_170_121 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_170_133 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_170_139 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_170_141 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_170_15 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_170_153 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_170_165 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_170_177 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_170_189 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_170_195 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_170_197 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_170_209 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_170_221 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_170_233 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_170_245 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_170_251 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_170_253 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_170_265 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_170_27 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_170_277 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_170_289 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_170_29 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_170_3 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_170_301 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_170_307 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_170_309 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_170_321 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_170_333 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_170_345 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_170_357 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_170_363 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_170_365 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_170_377 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_170_389 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_170_401 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_170_41 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_170_413 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_170_419 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_170_421 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_170_433 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_170_445 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_170_457 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_170_469 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_170_475 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_170_477 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_170_489 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_170_501 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_170_513 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_170_53 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_170_65 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_170_77 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_170_83 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_170_85 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_170_97 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_171_105 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_171_111 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_171_113 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_171_125 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_171_137 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_171_149 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_171_15 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_171_161 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_171_167 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_171_169 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_171_181 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_171_193 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_171_205 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_171_217 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_171_223 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_171_225 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_171_237 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_171_249 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_171_261 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_171_27 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_171_273 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_171_279 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_171_281 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_171_293 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_171_3 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_171_305 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_171_317 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_171_329 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_171_335 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_171_337 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_171_349 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_171_361 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_171_373 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_171_385 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_171_39 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_171_391 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_171_393 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_171_405 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_171_417 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_171_429 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_171_441 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_171_447 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_171_449 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_171_461 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_171_473 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_171_485 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_171_497 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_171_503 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_8 FILLER_171_505 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_4 FILLER_171_51 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_171_513 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_171_55 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_171_57 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_171_69 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_171_81 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_171_93 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_172_109 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_172_121 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_172_133 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_172_139 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_172_141 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_172_15 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_172_153 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_172_165 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_172_177 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_172_189 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_172_195 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_172_197 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_172_209 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_172_221 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_172_233 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_172_245 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_172_251 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_172_253 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_172_265 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_172_27 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_172_277 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_172_289 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_172_29 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_172_3 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_172_301 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_172_307 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_172_309 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_172_321 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_172_333 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_172_345 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_172_357 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_172_363 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_172_365 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_172_377 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_172_389 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_172_401 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_172_41 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_172_413 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_172_419 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_172_421 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_172_433 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_172_445 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_172_457 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_172_469 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_172_475 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_172_477 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_172_489 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_172_501 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_172_513 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_172_53 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_172_65 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_172_77 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_172_83 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_172_85 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_172_97 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_173_105 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_173_111 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_173_113 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_173_125 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_173_137 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_173_149 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_173_15 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_173_161 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_173_167 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_173_169 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_173_181 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_173_193 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_173_205 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_173_217 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_173_223 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_173_225 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_173_237 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_173_249 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_173_261 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_173_27 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_173_273 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_173_279 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_173_281 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_173_293 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_173_3 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_173_305 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_173_317 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_173_329 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_173_335 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_173_337 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_173_349 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_173_361 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_173_373 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_173_385 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_173_39 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_173_391 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_173_393 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_173_405 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_173_417 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_173_429 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_173_441 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_173_447 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_173_449 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_173_461 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_173_473 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_173_485 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_173_497 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_173_503 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_8 FILLER_173_505 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_4 FILLER_173_51 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_173_513 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_173_55 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_173_57 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_173_69 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_173_81 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_173_93 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_174_109 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_174_121 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_174_133 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_174_139 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_174_141 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_174_15 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_174_153 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_174_165 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_174_177 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_174_189 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_174_195 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_174_197 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_174_209 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_174_221 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_174_233 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_174_245 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_174_251 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_174_253 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_174_265 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_174_27 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_174_277 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_174_289 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_174_29 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_174_3 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_174_301 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_174_307 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_174_309 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_174_321 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_174_333 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_174_345 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_174_357 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_174_363 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_174_365 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_174_377 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_174_389 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_174_401 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_174_41 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_174_413 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_174_419 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_174_421 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_174_433 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_174_445 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_174_457 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_174_469 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_174_475 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_174_477 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_174_489 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_174_501 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_174_513 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_174_53 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_174_65 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_174_77 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_174_83 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_174_85 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_174_97 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_175_105 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_175_111 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_175_113 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_175_125 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_175_137 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_175_149 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_175_15 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_175_161 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_175_167 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_175_169 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_175_181 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_175_193 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_175_205 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_175_217 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_175_223 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_175_225 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_175_237 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_175_249 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_175_261 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_175_27 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_175_273 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_175_279 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_175_281 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_175_293 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_175_3 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_175_305 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_175_317 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_175_329 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_175_335 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_175_337 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_175_349 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_175_361 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_175_373 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_175_385 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_175_39 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_175_391 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_175_393 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_175_405 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_175_417 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_175_429 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_175_441 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_175_447 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_175_449 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_175_461 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_175_473 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_175_485 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_175_497 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_175_503 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_8 FILLER_175_505 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_4 FILLER_175_51 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_175_513 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_175_55 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_175_57 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_175_69 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_175_81 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_175_93 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_176_109 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_176_121 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_176_133 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_176_139 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_176_141 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_176_15 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_176_153 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_176_165 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_176_177 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_176_189 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_176_195 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_176_197 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_176_209 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_176_221 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_176_233 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_176_245 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_176_251 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_176_253 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_176_265 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_176_27 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_176_277 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_176_289 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_176_29 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_176_3 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_176_301 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_176_307 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_176_309 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_176_321 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_176_333 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_176_345 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_176_357 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_176_363 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_176_365 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_176_377 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_176_389 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_176_401 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_176_41 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_176_413 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_176_419 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_176_421 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_176_433 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_176_445 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_176_457 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_176_469 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_176_475 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_176_477 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_176_489 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_176_501 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_176_513 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_176_53 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_176_65 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_176_77 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_176_83 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_176_85 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_176_97 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_177_105 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_177_111 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_177_113 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_177_125 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_177_137 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_177_149 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_177_15 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_177_161 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_177_167 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_177_169 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_177_181 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_177_193 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_177_205 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_177_217 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_177_223 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_177_225 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_177_237 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_177_249 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_177_261 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_177_27 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_177_273 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_177_279 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_177_281 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_177_293 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_177_3 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_177_305 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_177_317 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_177_329 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_177_335 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_177_337 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_177_349 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_177_361 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_177_373 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_177_385 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_177_39 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_177_391 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_177_393 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_177_405 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_177_417 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_177_429 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_177_441 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_177_447 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_177_449 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_177_461 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_177_473 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_177_485 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_177_497 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_177_503 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_8 FILLER_177_505 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_4 FILLER_177_51 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_177_513 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_177_55 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_177_57 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_177_69 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_177_81 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_177_93 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_178_109 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_178_121 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_178_133 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_178_139 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_178_141 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_178_15 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_178_153 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_178_165 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_178_177 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_178_189 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_178_195 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_178_197 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_178_209 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_178_221 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_178_233 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_178_245 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_178_251 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_178_253 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_178_265 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_178_27 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_178_277 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_178_289 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_178_29 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_178_3 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_178_301 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_178_307 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_178_309 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_178_321 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_178_333 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_178_345 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_178_357 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_178_363 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_178_365 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_178_377 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_178_389 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_178_401 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_178_41 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_178_413 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_178_419 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_178_421 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_178_433 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_178_445 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_178_457 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_178_469 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_178_475 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_178_477 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_178_489 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_178_501 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_178_513 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_178_53 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_178_65 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_178_77 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_178_83 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_178_85 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_178_97 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_179_105 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_179_111 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_179_113 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_179_125 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_179_137 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_179_149 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_179_15 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_179_161 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_179_167 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_179_169 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_179_181 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_179_193 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_179_205 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_179_217 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_179_223 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_179_225 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_179_237 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_179_249 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_179_261 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_179_27 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_179_273 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_179_279 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_179_281 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_179_293 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_179_3 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_179_305 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_179_317 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_179_329 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_179_335 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_179_337 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_179_349 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_179_361 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_179_373 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_179_385 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_179_39 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_179_391 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_179_393 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_179_405 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_179_417 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_179_429 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_179_441 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_179_447 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_179_449 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_179_461 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_179_473 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_179_485 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_179_497 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_179_503 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_8 FILLER_179_505 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_4 FILLER_179_51 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_179_513 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_179_55 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_179_57 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_179_69 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_179_81 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_179_93 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_17_105 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_17_111 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_17_113 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_17_125 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_17_137 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_17_149 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_17_15 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_17_161 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_17_167 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_17_169 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_17_181 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_17_193 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_17_205 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_17_217 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_17_223 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_17_225 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_17_237 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_17_249 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_17_261 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_17_27 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_17_273 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_17_279 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_17_281 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_17_293 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_17_3 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_17_305 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_17_317 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_17_329 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_17_335 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_17_337 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_17_349 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_17_361 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_17_373 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_17_385 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_17_39 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_17_391 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_17_393 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_17_405 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_17_417 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_17_429 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_17_441 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_17_447 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_17_449 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_17_461 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_17_473 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_17_485 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_17_497 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_17_503 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_8 FILLER_17_505 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_4 FILLER_17_51 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_17_513 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_17_55 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_17_57 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_17_69 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_17_81 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_17_93 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_180_109 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_180_121 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_180_133 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_180_139 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_180_141 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_180_15 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_180_153 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_180_165 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_180_177 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_180_189 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_180_195 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_180_197 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_180_209 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_180_221 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_180_233 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_180_245 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_180_251 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_180_253 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_180_265 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_180_27 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_180_277 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_180_289 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_180_29 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_180_3 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_180_301 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_180_307 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_180_309 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_180_321 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_180_333 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_180_345 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_180_357 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_180_363 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_180_365 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_180_377 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_180_389 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_180_401 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_180_41 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_180_413 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_180_419 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_180_421 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_180_433 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_180_445 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_180_457 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_180_469 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_180_475 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_180_477 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_180_489 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_180_501 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_180_513 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_180_53 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_180_65 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_180_77 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_180_83 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_180_85 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_180_97 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_181_105 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_181_111 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_181_113 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_181_125 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_181_137 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_181_149 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_181_15 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_181_161 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_181_167 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_181_169 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_181_181 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_181_193 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_181_205 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_181_217 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_181_223 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_181_225 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_181_237 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_181_249 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_181_261 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_181_27 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_181_273 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_181_279 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_181_281 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_181_293 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_181_3 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_181_305 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_181_317 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_181_329 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_181_335 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_181_337 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_181_349 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_181_361 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_181_373 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_181_385 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_181_39 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_181_391 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_181_393 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_181_405 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_181_417 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_181_429 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_181_441 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_181_447 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_181_449 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_181_461 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_181_473 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_181_485 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_181_497 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_181_503 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_8 FILLER_181_505 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_4 FILLER_181_51 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_181_513 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_181_55 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_181_57 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_181_69 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_181_81 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_181_93 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_182_109 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_182_121 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_182_133 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_182_139 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_182_141 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_182_15 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_182_153 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_182_165 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_182_177 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_182_189 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_182_195 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_182_197 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_182_209 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_182_221 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_182_233 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_182_245 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_182_251 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_182_253 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_182_265 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_182_27 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_182_277 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_182_289 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_182_29 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_182_3 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_182_301 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_182_307 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_182_309 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_182_321 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_182_333 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_182_345 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_182_357 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_182_363 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_182_365 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_182_377 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_182_389 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_182_401 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_182_41 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_182_413 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_182_419 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_182_421 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_182_433 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_182_445 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_182_457 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_182_469 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_182_475 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_182_477 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_182_489 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_182_501 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_182_513 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_182_53 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_182_65 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_182_77 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_182_83 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_182_85 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_182_97 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_183_105 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_183_111 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_183_113 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_183_125 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_183_137 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_183_149 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_183_15 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_183_161 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_183_167 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_183_169 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_183_181 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_183_193 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_183_205 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_183_217 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_183_223 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_183_225 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_183_237 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_183_249 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_183_261 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_183_27 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_183_273 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_183_279 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_183_281 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_183_293 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_183_3 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_183_305 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_183_317 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_183_329 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_183_335 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_183_337 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_183_349 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_183_361 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_183_373 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_183_385 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_183_39 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_183_391 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_183_393 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_183_405 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_183_417 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_183_429 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_183_441 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_183_447 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_183_449 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_183_461 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_183_473 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_183_485 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_183_497 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_183_503 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_8 FILLER_183_505 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_4 FILLER_183_51 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_183_513 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_183_55 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_183_57 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_183_69 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_183_81 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_183_93 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_184_109 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_184_121 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_184_133 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_184_139 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_184_141 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_184_15 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_184_153 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_184_165 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_184_177 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_184_189 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_184_195 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_184_197 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_184_209 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_184_221 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_184_233 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_184_245 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_184_251 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_184_253 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_184_265 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_184_27 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_184_277 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_184_289 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_184_29 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_184_3 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_184_301 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_184_307 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_184_309 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_184_321 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_184_333 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_184_345 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_184_357 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_184_363 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_184_365 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_184_377 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_184_389 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_184_401 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_184_41 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_184_413 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_184_419 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_184_421 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_184_433 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_184_445 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_184_457 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_184_469 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_184_475 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_184_477 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_184_489 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_184_501 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_184_513 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_184_53 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_184_65 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_184_77 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_184_83 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_184_85 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_184_97 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_185_105 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_185_111 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_185_113 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_185_125 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_185_137 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_185_149 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_185_15 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_185_161 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_185_167 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_185_169 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_185_181 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_185_193 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_185_205 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_185_217 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_185_223 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_185_225 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_185_237 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_185_249 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_185_261 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_185_27 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_185_273 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_185_279 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_185_281 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_185_293 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_185_3 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_185_305 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_185_317 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_185_329 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_185_335 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_185_337 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_185_349 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_185_361 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_185_373 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_185_385 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_185_39 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_185_391 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_185_393 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_185_405 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_185_417 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_185_429 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_185_441 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_185_447 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_185_449 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_185_461 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_185_473 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_185_485 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_185_497 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_185_503 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_8 FILLER_185_505 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_4 FILLER_185_51 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_185_513 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_185_55 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_185_57 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_185_69 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_185_81 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_185_93 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_186_109 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_186_121 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_186_133 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_186_139 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_186_141 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_186_15 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_186_153 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_186_165 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_186_177 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_186_189 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_186_195 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_186_197 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_186_209 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_186_221 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_186_233 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_186_245 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_186_251 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_186_253 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_186_265 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_186_27 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_186_277 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_186_289 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_186_29 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_186_3 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_186_301 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_186_307 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_186_309 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_186_321 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_186_333 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_186_345 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_186_357 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_186_363 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_186_365 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_186_377 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_186_389 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_186_401 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_186_41 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_186_413 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_186_419 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_186_421 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_186_433 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_186_445 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_186_457 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_186_469 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_186_475 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_186_477 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_186_489 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_186_501 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_186_513 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_186_53 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_186_65 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_186_77 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_186_83 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_186_85 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_186_97 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_187_105 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_187_111 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_187_113 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_4 FILLER_187_125 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_4 FILLER_187_149 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_187_15 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_187_155 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_187_167 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_8 FILLER_187_169 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_187_177 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_4 FILLER_187_182 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_187_206 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_187_218 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_187_225 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_187_237 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_187_249 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_187_261 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_187_27 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_187_273 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_187_279 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_187_281 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_187_293 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_187_3 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_187_305 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_187_317 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_187_329 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_187_335 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_187_337 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_187_349 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_187_361 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_187_373 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_187_385 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_187_39 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_187_391 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_187_393 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_187_405 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_187_417 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_187_429 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_187_441 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_187_447 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_187_449 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_187_461 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_187_473 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_187_485 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_187_497 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_187_503 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_8 FILLER_187_505 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_4 FILLER_187_51 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_187_513 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_187_55 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_187_57 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_187_69 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_187_81 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_187_93 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_188_109 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_188_121 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_188_133 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_188_139 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_188_141 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_188_15 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_188_153 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_8 FILLER_188_165 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_188_173 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_188_176 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_8 FILLER_188_188 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_188_197 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_188_209 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_188_221 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_2 FILLER_188_233 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_188_237 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_188_249 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_188_253 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_188_265 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_188_27 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_188_277 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_8 FILLER_188_289 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_188_29 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_2 FILLER_188_297 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_188_3 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_188_301 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_188_307 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_188_309 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_188_321 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_188_333 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_188_345 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_188_357 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_188_363 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_188_365 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_188_377 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_188_389 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_188_401 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_188_41 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_188_413 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_188_419 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_188_421 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_188_433 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_188_445 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_188_457 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_188_469 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_188_475 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_188_477 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_188_489 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_188_501 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_188_513 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_8 FILLER_188_53 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_188_61 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_188_64 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_8 FILLER_188_76 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_188_85 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_188_97 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_8 FILLER_189_102 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_2 FILLER_189_110 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_189_113 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_189_125 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_189_137 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_189_149 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_189_15 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_189_161 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_189_167 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_2 FILLER_189_169 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_189_188 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_189_200 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_189_212 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_189_225 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_4 FILLER_189_230 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_189_251 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_189_263 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_189_27 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_4 FILLER_189_275 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_189_279 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_8 FILLER_189_281 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_189_289 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_4 FILLER_189_292 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_189_3 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_189_313 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_8 FILLER_189_325 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_189_333 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_189_337 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_189_349 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_189_361 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_189_373 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_189_385 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_189_39 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_189_391 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_189_393 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_189_405 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_189_417 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_189_429 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_189_441 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_189_447 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_189_449 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_189_461 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_189_473 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_189_485 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_189_497 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_189_503 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_8 FILLER_189_505 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_4 FILLER_189_51 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_189_513 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_189_55 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_4 FILLER_189_57 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_189_78 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_189_90 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_18_109 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_18_121 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_18_133 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_18_139 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_18_141 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_18_15 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_18_153 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_18_165 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_18_177 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_18_189 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_18_195 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_18_197 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_18_209 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_18_221 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_18_233 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_18_245 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_18_251 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_18_253 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_18_265 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_18_27 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_18_277 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_18_289 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_18_29 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_18_3 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_18_301 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_18_307 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_18_309 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_18_321 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_18_333 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_18_345 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_18_357 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_18_363 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_18_365 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_18_377 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_18_389 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_18_401 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_18_41 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_18_413 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_18_419 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_18_421 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_18_433 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_18_445 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_18_457 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_18_469 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_18_475 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_18_477 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_18_489 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_18_501 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_18_513 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_18_53 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_18_65 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_18_77 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_18_83 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_18_85 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_18_97 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_190_109 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_190_121 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_190_133 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_190_139 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_190_141 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_190_15 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_190_153 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_190_165 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_4 FILLER_190_170 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_2 FILLER_190_194 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_190_197 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_190_209 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_190_221 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_190_233 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_190_245 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_190_251 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_190_253 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_190_265 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_190_27 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_190_277 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_190_289 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_190_29 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_190_3 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_190_301 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_190_307 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_190_309 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_190_321 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_190_333 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_190_345 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_190_357 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_190_363 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_190_365 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_190_377 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_190_389 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_190_401 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_190_41 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_190_413 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_190_419 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_190_421 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_190_433 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_190_445 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_190_457 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_190_469 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_190_475 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_190_477 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_190_489 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_190_501 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_190_513 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_190_53 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_190_61 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_8 FILLER_190_73 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_190_81 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_190_85 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_190_97 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_191_105 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_191_111 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_191_113 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_191_125 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_191_137 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_191_149 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_191_15 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_191_161 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_191_167 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_191_169 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_191_177 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_191_189 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_191_201 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_8 FILLER_191_213 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_191_221 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_191_225 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_191_237 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_191_249 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_191_261 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_191_27 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_191_273 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_191_279 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_191_281 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_191_293 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_191_3 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_191_305 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_191_317 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_191_329 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_191_335 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_191_337 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_191_349 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_191_361 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_191_373 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_191_385 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_191_39 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_191_391 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_191_393 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_191_405 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_191_417 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_191_429 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_191_441 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_191_447 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_191_449 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_191_461 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_191_473 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_191_485 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_191_497 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_191_503 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_8 FILLER_191_505 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_4 FILLER_191_51 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_191_513 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_191_55 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_191_57 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_191_69 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_191_81 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_191_93 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_192_109 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_192_121 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_192_133 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_192_139 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_192_141 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_192_15 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_192_153 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_192_165 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_192_177 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_192_189 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_192_195 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_192_197 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_192_209 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_192_221 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_192_233 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_192_245 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_192_251 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_192_253 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_192_265 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_192_27 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_192_277 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_192_289 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_192_29 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_192_3 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_192_301 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_192_307 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_192_309 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_192_321 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_192_333 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_192_345 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_192_357 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_192_363 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_192_365 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_192_377 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_192_389 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_192_401 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_192_41 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_192_413 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_192_419 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_192_421 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_192_433 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_192_445 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_192_457 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_192_469 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_192_475 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_192_477 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_192_489 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_192_501 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_192_513 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_192_53 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_192_65 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_192_77 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_192_83 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_192_85 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_192_97 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_193_109 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_193_113 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_193_125 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_193_137 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_193_141 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_193_15 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_193_153 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_193_165 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_193_169 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_193_181 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_193_193 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_193_197 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_193_209 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_193_221 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_193_225 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_193_237 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_193_249 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_193_253 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_193_265 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_193_27 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_193_277 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_193_281 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_193_29 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_193_293 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_193_3 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_193_305 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_193_309 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_193_321 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_193_333 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_193_337 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_193_349 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_193_361 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_193_365 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_193_377 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_193_389 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_193_393 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_193_405 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_193_41 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_193_417 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_193_421 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_193_433 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_193_445 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_193_449 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_193_461 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_193_473 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_193_477 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_193_489 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_193_501 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_8 FILLER_193_505 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_193_513 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_193_53 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_193_57 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_193_69 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_193_81 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_193_85 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_193_97 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_19_105 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_19_111 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_19_113 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_19_125 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_19_137 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_19_149 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_19_15 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_19_161 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_19_167 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_19_169 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_19_181 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_19_193 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_19_205 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_19_217 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_19_223 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_19_225 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_19_237 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_19_249 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_19_261 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_19_27 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_19_273 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_19_279 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_19_281 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_19_293 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_19_3 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_19_305 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_19_317 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_19_329 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_19_335 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_19_337 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_19_349 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_19_361 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_19_373 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_19_385 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_19_39 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_19_391 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_19_393 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_19_405 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_19_417 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_19_429 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_19_441 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_19_447 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_19_449 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_19_461 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_19_473 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_19_485 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_19_497 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_19_503 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_8 FILLER_19_505 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_4 FILLER_19_51 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_19_513 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_19_55 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_19_57 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_19_69 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_19_81 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_19_93 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_1_105 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_1_111 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_1_113 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_1_125 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_1_137 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_1_149 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_1_15 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_1_161 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_1_167 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_1_169 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_1_181 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_1_193 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_1_205 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_1_217 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_1_223 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_1_225 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_1_237 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_1_249 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_1_261 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_1_27 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_1_273 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_1_279 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_1_281 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_1_293 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_1_3 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_1_305 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_1_317 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_1_329 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_1_335 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_1_337 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_1_349 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_1_361 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_1_373 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_1_385 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_1_39 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_1_391 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_1_393 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_1_405 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_1_417 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_1_429 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_1_441 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_1_447 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_1_449 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_1_461 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_1_473 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_1_485 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_1_497 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_1_503 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_8 FILLER_1_505 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_4 FILLER_1_51 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_1_513 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_1_55 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_1_57 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_1_69 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_1_81 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_1_93 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_20_109 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_20_121 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_20_133 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_20_139 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_20_141 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_20_15 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_20_153 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_20_165 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_20_177 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_20_189 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_20_195 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_20_197 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_20_209 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_20_221 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_20_233 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_20_245 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_20_251 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_20_253 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_20_265 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_20_27 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_20_277 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_20_289 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_20_29 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_20_3 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_20_301 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_20_307 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_20_309 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_20_321 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_20_333 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_20_345 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_20_357 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_20_363 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_20_365 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_20_377 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_20_389 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_20_401 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_20_41 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_20_413 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_20_419 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_20_421 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_20_433 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_20_445 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_20_457 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_20_469 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_20_475 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_20_477 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_20_489 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_20_501 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_20_513 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_20_53 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_20_65 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_20_77 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_20_83 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_20_85 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_20_97 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_21_105 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_21_111 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_21_113 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_21_125 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_21_137 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_21_149 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_21_15 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_21_161 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_21_167 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_21_169 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_21_181 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_21_193 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_21_205 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_21_217 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_21_223 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_21_225 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_21_237 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_21_249 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_21_261 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_21_27 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_21_273 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_21_279 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_21_281 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_21_293 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_21_3 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_21_305 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_21_317 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_21_329 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_21_335 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_21_337 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_21_349 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_21_361 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_21_373 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_21_385 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_21_39 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_21_391 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_21_393 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_21_405 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_21_417 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_21_429 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_21_441 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_21_447 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_21_449 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_21_461 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_21_473 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_21_485 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_21_497 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_21_503 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_8 FILLER_21_505 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_4 FILLER_21_51 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_21_513 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_21_55 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_21_57 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_21_69 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_21_81 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_21_93 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_22_109 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_22_121 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_22_133 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_22_139 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_22_141 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_22_15 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_22_153 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_22_165 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_22_177 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_22_189 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_22_195 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_22_197 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_22_209 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_22_221 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_22_233 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_22_245 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_22_251 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_22_253 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_22_265 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_22_27 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_22_277 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_22_289 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_22_29 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_22_3 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_22_301 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_22_307 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_22_309 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_22_321 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_22_333 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_22_345 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_22_357 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_22_363 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_22_365 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_22_377 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_22_389 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_22_401 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_22_41 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_22_413 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_22_419 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_22_421 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_22_433 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_22_445 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_22_457 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_22_469 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_22_475 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_22_477 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_22_489 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_22_501 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_22_513 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_22_53 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_22_65 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_22_77 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_22_83 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_22_85 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_22_97 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_23_105 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_23_111 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_23_113 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_23_125 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_23_137 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_23_149 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_23_15 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_23_161 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_23_167 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_23_169 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_23_181 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_23_193 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_23_205 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_23_217 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_23_223 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_23_225 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_23_237 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_23_249 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_23_261 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_23_27 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_23_273 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_23_279 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_23_281 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_23_293 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_23_3 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_23_305 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_23_317 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_23_329 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_23_335 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_23_337 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_23_349 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_23_361 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_23_373 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_23_385 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_23_39 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_23_391 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_23_393 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_23_405 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_23_417 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_23_429 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_23_441 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_23_447 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_23_449 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_23_461 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_23_473 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_23_485 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_23_497 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_23_503 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_8 FILLER_23_505 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_4 FILLER_23_51 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_23_513 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_23_55 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_23_57 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_23_69 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_23_81 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_23_93 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_24_109 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_24_121 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_24_133 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_24_139 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_24_141 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_24_15 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_24_153 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_24_165 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_24_177 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_24_189 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_24_195 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_24_197 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_24_209 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_24_221 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_24_233 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_24_245 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_24_251 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_24_253 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_24_265 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_24_27 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_24_277 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_24_289 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_24_29 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_24_3 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_24_301 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_24_307 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_24_309 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_24_321 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_24_333 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_24_345 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_24_357 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_24_363 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_24_365 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_24_377 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_24_389 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_24_401 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_24_41 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_24_413 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_24_419 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_24_421 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_24_433 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_24_445 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_24_457 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_24_469 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_24_475 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_24_477 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_24_489 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_24_501 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_24_513 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_24_53 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_24_65 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_24_77 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_24_83 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_24_85 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_24_97 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_25_105 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_25_111 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_25_113 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_25_125 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_25_137 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_25_149 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_25_15 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_25_161 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_25_167 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_25_169 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_25_181 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_25_193 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_25_205 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_25_217 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_25_223 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_25_225 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_25_237 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_25_249 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_25_261 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_25_27 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_25_273 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_25_279 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_25_281 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_25_293 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_25_3 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_25_305 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_25_317 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_25_329 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_25_335 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_25_337 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_25_349 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_25_361 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_25_373 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_25_385 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_25_39 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_25_391 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_25_393 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_25_405 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_25_417 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_25_429 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_25_441 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_25_447 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_25_449 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_25_461 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_25_473 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_25_485 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_25_497 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_25_503 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_8 FILLER_25_505 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_4 FILLER_25_51 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_25_513 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_25_55 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_25_57 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_25_69 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_25_81 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_25_93 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_26_109 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_26_121 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_26_133 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_26_139 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_26_141 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_26_15 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_26_153 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_26_165 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_26_177 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_26_189 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_26_195 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_26_197 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_26_209 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_26_221 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_26_233 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_26_245 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_26_251 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_26_253 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_26_265 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_26_27 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_26_277 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_26_289 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_26_29 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_26_3 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_26_301 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_26_307 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_26_309 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_26_321 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_26_333 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_26_345 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_26_357 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_26_363 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_26_365 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_26_377 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_26_389 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_26_401 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_26_41 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_26_413 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_26_419 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_26_421 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_26_433 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_26_445 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_26_457 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_26_469 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_26_475 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_26_477 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_26_489 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_26_501 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_26_513 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_26_53 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_26_65 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_26_77 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_26_83 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_26_85 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_26_97 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_27_105 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_27_111 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_27_113 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_27_125 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_27_137 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_27_149 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_27_15 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_27_161 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_27_167 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_27_169 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_27_181 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_27_193 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_27_205 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_27_217 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_27_223 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_27_225 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_27_237 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_27_249 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_27_261 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_27_27 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_27_273 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_27_279 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_27_281 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_27_293 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_27_3 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_27_305 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_27_317 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_27_329 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_27_335 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_27_337 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_27_349 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_27_361 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_27_373 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_27_385 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_27_39 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_27_391 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_27_393 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_27_405 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_27_417 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_27_429 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_27_441 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_27_447 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_27_449 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_27_461 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_27_473 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_27_485 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_27_497 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_27_503 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_8 FILLER_27_505 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_4 FILLER_27_51 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_27_513 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_27_55 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_27_57 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_27_69 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_27_81 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_27_93 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_28_109 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_28_121 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_28_133 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_28_139 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_28_141 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_28_15 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_28_153 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_28_165 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_28_177 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_28_189 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_28_195 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_28_197 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_28_209 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_28_221 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_28_233 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_28_245 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_28_251 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_28_253 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_28_265 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_28_27 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_28_277 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_28_289 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_28_29 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_28_3 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_28_301 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_28_307 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_28_309 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_28_321 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_28_333 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_28_345 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_28_357 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_28_363 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_28_365 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_28_377 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_28_389 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_28_401 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_28_41 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_28_413 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_28_419 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_28_421 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_28_433 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_28_445 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_28_457 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_28_469 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_28_475 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_28_477 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_28_489 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_28_501 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_28_513 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_28_53 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_28_65 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_28_77 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_28_83 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_28_85 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_28_97 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_29_105 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_29_111 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_29_113 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_29_125 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_29_137 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_29_149 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_29_15 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_29_161 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_29_167 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_29_169 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_29_181 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_29_193 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_29_205 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_29_217 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_29_223 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_29_225 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_29_237 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_29_249 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_29_261 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_29_27 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_29_273 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_29_279 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_29_281 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_29_293 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_29_3 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_29_305 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_29_317 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_29_329 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_29_335 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_29_337 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_29_349 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_29_361 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_29_373 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_29_385 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_29_39 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_29_391 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_29_393 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_29_405 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_29_417 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_29_429 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_29_441 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_29_447 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_29_449 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_29_461 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_29_473 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_29_485 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_29_497 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_29_503 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_8 FILLER_29_505 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_4 FILLER_29_51 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_29_513 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_29_55 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_29_57 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_29_69 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_29_81 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_29_93 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_2_109 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_2_121 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_2_133 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_2_139 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_2_141 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_2_15 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_2_153 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_2_165 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_2_177 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_2_189 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_2_195 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_2_197 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_2_209 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_2_221 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_2_233 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_2_245 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_2_251 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_2_253 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_2_265 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_2_27 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_2_277 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_2_289 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_2_29 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_2_3 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_2_301 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_2_307 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_2_309 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_2_321 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_2_333 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_2_345 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_2_357 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_2_363 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_2_365 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_2_377 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_2_389 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_2_401 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_2_41 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_2_413 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_2_419 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_2_421 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_2_433 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_2_445 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_2_457 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_2_469 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_2_475 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_2_477 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_2_489 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_2_501 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_2_513 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_2_53 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_2_65 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_2_77 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_2_83 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_2_85 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_2_97 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_30_109 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_30_121 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_30_133 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_30_139 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_30_141 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_30_15 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_30_153 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_30_165 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_30_177 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_30_189 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_30_195 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_30_197 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_30_209 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_30_221 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_30_233 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_30_245 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_30_251 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_30_253 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_30_265 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_30_27 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_30_277 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_30_289 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_30_29 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_30_3 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_30_301 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_30_307 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_30_309 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_30_321 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_30_333 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_30_345 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_30_357 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_30_363 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_30_365 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_30_377 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_30_389 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_30_401 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_30_41 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_30_413 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_30_419 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_30_421 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_30_433 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_30_445 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_30_457 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_30_469 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_30_475 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_30_477 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_30_489 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_30_501 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_30_513 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_30_53 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_30_65 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_30_77 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_30_83 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_30_85 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_30_97 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_31_105 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_31_111 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_31_113 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_31_125 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_31_137 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_31_149 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_31_15 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_31_161 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_31_167 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_31_169 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_31_181 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_31_193 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_31_205 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_31_217 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_31_223 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_31_225 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_31_237 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_31_249 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_31_261 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_31_27 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_31_273 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_31_279 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_31_281 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_31_293 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_31_3 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_31_305 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_31_317 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_31_329 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_31_335 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_31_337 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_31_349 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_31_361 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_31_373 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_31_385 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_31_39 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_31_391 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_31_393 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_31_405 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_31_417 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_31_429 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_31_441 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_31_447 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_31_449 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_31_461 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_31_473 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_31_485 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_31_497 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_31_503 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_8 FILLER_31_505 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_4 FILLER_31_51 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_31_513 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_31_55 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_31_57 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_31_69 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_31_81 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_31_93 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_32_109 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_32_121 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_32_133 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_32_139 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_32_141 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_32_15 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_32_153 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_32_165 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_32_177 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_32_189 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_32_195 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_32_197 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_32_209 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_32_221 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_32_233 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_32_245 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_32_251 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_32_253 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_32_265 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_32_27 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_32_277 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_32_289 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_32_29 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_32_3 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_32_301 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_32_307 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_32_309 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_32_321 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_32_333 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_32_345 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_32_357 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_32_363 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_32_365 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_32_377 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_32_389 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_32_401 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_32_41 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_32_413 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_32_419 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_32_421 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_32_433 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_32_445 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_32_457 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_32_469 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_32_475 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_32_477 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_32_489 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_32_501 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_32_513 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_32_53 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_32_65 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_32_77 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_32_83 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_32_85 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_32_97 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_33_105 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_33_111 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_33_113 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_33_125 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_33_137 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_33_149 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_33_15 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_33_161 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_33_167 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_33_169 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_33_181 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_33_193 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_33_205 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_33_217 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_33_223 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_33_225 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_33_237 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_33_249 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_33_261 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_33_27 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_33_273 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_33_279 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_33_281 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_33_293 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_33_3 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_33_305 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_33_317 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_33_329 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_33_335 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_33_337 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_33_349 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_33_361 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_33_373 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_33_385 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_33_39 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_33_391 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_33_393 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_33_405 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_33_417 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_33_429 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_33_441 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_33_447 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_33_449 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_33_461 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_33_473 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_33_485 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_33_497 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_33_503 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_8 FILLER_33_505 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_4 FILLER_33_51 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_33_513 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_33_55 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_33_57 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_33_69 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_33_81 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_33_93 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_34_109 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_34_121 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_34_133 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_34_139 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_34_141 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_34_15 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_34_153 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_34_165 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_34_177 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_34_189 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_34_195 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_34_197 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_34_209 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_34_221 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_34_233 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_34_245 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_34_251 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_34_253 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_34_265 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_34_27 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_34_277 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_34_289 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_34_29 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_34_3 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_34_301 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_34_307 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_34_309 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_34_321 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_34_333 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_34_345 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_34_357 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_34_363 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_34_365 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_34_377 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_34_389 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_34_401 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_34_41 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_34_413 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_34_419 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_34_421 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_34_433 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_34_445 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_34_457 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_34_469 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_34_475 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_34_477 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_34_489 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_34_501 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_34_513 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_34_53 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_34_65 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_34_77 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_34_83 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_34_85 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_34_97 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_35_105 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_35_111 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_35_113 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_35_125 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_35_137 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_35_149 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_35_15 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_35_161 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_35_167 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_35_169 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_35_181 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_35_193 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_35_205 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_35_217 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_35_223 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_35_225 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_35_237 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_35_249 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_35_261 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_35_27 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_35_273 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_35_279 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_35_281 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_35_293 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_35_3 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_35_305 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_35_317 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_35_329 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_35_335 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_35_337 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_35_349 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_35_361 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_35_373 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_35_385 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_35_39 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_35_391 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_35_393 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_35_405 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_35_417 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_35_429 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_35_441 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_35_447 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_35_449 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_35_461 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_35_473 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_35_485 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_35_497 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_35_503 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_8 FILLER_35_505 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_4 FILLER_35_51 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_35_513 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_35_55 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_35_57 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_35_69 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_35_81 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_35_93 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_36_109 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_36_121 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_36_133 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_36_139 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_36_141 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_36_15 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_36_153 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_36_165 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_36_177 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_36_189 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_36_195 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_36_197 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_36_209 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_36_221 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_36_233 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_36_245 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_36_251 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_36_253 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_36_265 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_36_27 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_36_277 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_36_289 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_36_29 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_36_3 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_36_301 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_36_307 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_36_309 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_36_321 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_36_333 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_36_345 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_36_357 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_36_363 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_36_365 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_36_377 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_36_389 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_36_401 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_36_41 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_36_413 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_36_419 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_36_421 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_36_433 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_36_445 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_36_457 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_36_469 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_36_475 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_36_477 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_36_489 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_36_501 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_36_513 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_36_53 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_36_65 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_36_77 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_36_83 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_36_85 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_36_97 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_37_105 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_37_111 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_37_113 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_37_125 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_37_137 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_37_149 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_37_15 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_37_161 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_37_167 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_37_169 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_37_181 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_37_193 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_37_205 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_37_217 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_37_223 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_37_225 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_37_237 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_37_249 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_37_261 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_37_27 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_37_273 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_37_279 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_37_281 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_37_293 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_37_3 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_37_305 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_37_317 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_37_329 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_37_335 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_37_337 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_37_349 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_37_361 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_37_373 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_37_385 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_37_39 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_37_391 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_37_393 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_37_405 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_37_417 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_37_429 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_37_441 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_37_447 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_37_449 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_37_461 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_37_473 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_37_485 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_37_497 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_37_503 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_8 FILLER_37_505 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_4 FILLER_37_51 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_37_513 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_37_55 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_37_57 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_37_69 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_37_81 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_37_93 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_38_109 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_38_121 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_38_133 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_38_139 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_38_141 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_38_15 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_38_153 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_38_165 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_38_177 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_38_189 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_38_195 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_38_197 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_38_209 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_38_221 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_38_233 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_38_245 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_38_251 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_38_253 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_38_265 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_38_27 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_38_277 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_38_289 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_38_29 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_38_3 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_38_301 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_38_307 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_38_309 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_38_321 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_38_333 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_38_345 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_38_357 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_38_363 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_38_365 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_38_377 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_38_389 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_38_401 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_38_41 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_38_413 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_38_419 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_38_421 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_38_433 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_38_445 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_38_457 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_38_469 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_38_475 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_38_477 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_38_489 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_38_501 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_38_513 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_38_53 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_38_65 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_38_77 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_38_83 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_38_85 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_38_97 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_39_105 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_39_111 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_39_113 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_39_125 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_39_137 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_39_149 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_39_15 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_39_161 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_39_167 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_39_169 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_39_181 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_39_193 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_39_205 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_39_217 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_39_223 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_39_225 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_39_237 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_39_249 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_39_261 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_39_27 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_39_273 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_39_279 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_39_281 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_39_293 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_39_3 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_39_305 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_39_317 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_39_329 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_39_335 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_39_337 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_39_349 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_39_361 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_39_373 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_39_385 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_39_39 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_39_391 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_39_393 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_39_405 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_39_417 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_39_429 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_39_441 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_39_447 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_39_449 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_39_461 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_39_473 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_39_485 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_39_497 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_39_503 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_8 FILLER_39_505 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_4 FILLER_39_51 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_39_513 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_39_55 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_39_57 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_39_69 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_39_81 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_39_93 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_3_105 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_3_111 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_3_113 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_3_125 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_3_137 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_3_149 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_3_15 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_3_161 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_3_167 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_3_169 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_3_181 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_3_193 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_3_205 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_3_217 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_3_223 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_3_225 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_3_237 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_3_249 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_3_261 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_3_27 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_3_273 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_3_279 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_3_281 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_3_293 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_3_3 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_3_305 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_3_317 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_3_329 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_3_335 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_3_337 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_3_349 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_3_361 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_3_373 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_3_385 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_3_39 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_3_391 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_3_393 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_3_405 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_3_417 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_3_429 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_3_441 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_3_447 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_3_449 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_3_461 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_3_473 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_3_485 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_3_497 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_3_503 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_8 FILLER_3_505 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_4 FILLER_3_51 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_3_513 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_3_55 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_3_57 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_3_69 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_3_81 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_3_93 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_40_109 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_40_121 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_40_133 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_40_139 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_40_141 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_40_15 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_40_153 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_40_165 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_40_177 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_40_189 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_40_195 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_40_197 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_40_209 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_40_221 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_40_233 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_40_245 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_40_251 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_40_253 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_40_265 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_40_27 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_40_277 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_40_289 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_40_29 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_40_3 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_40_301 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_40_307 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_40_309 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_40_321 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_40_333 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_40_345 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_40_357 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_40_363 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_40_365 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_40_377 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_40_389 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_40_401 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_40_41 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_40_413 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_40_419 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_40_421 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_40_433 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_40_445 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_40_457 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_40_469 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_40_475 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_40_477 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_40_489 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_40_501 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_40_513 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_40_53 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_40_65 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_40_77 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_40_83 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_40_85 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_40_97 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_41_105 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_41_111 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_41_113 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_41_125 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_41_137 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_41_149 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_41_15 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_41_161 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_41_167 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_41_169 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_41_181 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_41_193 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_41_205 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_41_217 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_41_223 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_41_225 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_41_237 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_41_249 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_41_261 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_41_27 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_41_273 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_41_279 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_41_281 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_41_293 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_41_3 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_41_305 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_41_317 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_41_329 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_41_335 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_41_337 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_41_349 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_41_361 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_41_373 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_41_385 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_41_39 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_41_391 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_41_393 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_41_405 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_41_417 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_41_429 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_41_441 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_41_447 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_41_449 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_41_461 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_41_473 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_41_485 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_41_497 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_41_503 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_8 FILLER_41_505 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_4 FILLER_41_51 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_41_513 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_41_55 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_41_57 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_41_69 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_41_81 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_41_93 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_42_109 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_42_121 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_42_133 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_42_139 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_42_141 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_42_15 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_42_153 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_42_165 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_42_177 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_42_189 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_42_195 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_42_197 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_42_209 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_42_221 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_42_233 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_42_245 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_42_251 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_42_253 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_42_265 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_42_27 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_42_277 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_42_289 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_42_29 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_42_3 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_42_301 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_42_307 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_42_309 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_42_321 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_42_333 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_42_345 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_42_357 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_42_363 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_42_365 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_42_377 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_42_389 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_42_401 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_42_41 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_42_413 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_42_419 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_42_421 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_42_433 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_42_445 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_42_457 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_42_469 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_42_475 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_42_477 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_42_489 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_42_501 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_42_513 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_42_53 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_42_65 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_42_77 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_42_83 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_42_85 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_42_97 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_43_105 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_43_111 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_43_113 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_43_125 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_43_137 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_43_149 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_43_15 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_43_161 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_43_167 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_43_169 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_43_181 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_43_193 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_43_205 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_43_217 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_43_223 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_43_225 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_43_237 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_43_249 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_43_261 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_43_27 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_43_273 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_43_279 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_43_281 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_43_293 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_43_3 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_43_305 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_43_317 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_43_329 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_43_335 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_43_337 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_43_349 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_43_361 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_43_373 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_43_385 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_43_39 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_43_391 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_43_393 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_43_405 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_43_417 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_43_429 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_43_441 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_43_447 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_43_449 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_43_461 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_43_473 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_43_485 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_43_497 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_43_503 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_8 FILLER_43_505 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_4 FILLER_43_51 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_43_513 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_43_55 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_43_57 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_43_69 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_43_81 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_43_93 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_44_109 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_44_121 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_44_133 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_44_139 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_44_141 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_44_15 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_44_153 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_44_165 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_44_177 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_44_189 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_44_195 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_44_197 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_44_209 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_44_221 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_44_233 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_44_245 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_44_251 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_44_253 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_44_265 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_44_27 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_44_277 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_44_289 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_44_29 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_44_3 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_44_301 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_44_307 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_44_309 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_44_321 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_44_333 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_44_345 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_44_357 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_44_363 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_44_365 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_44_377 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_44_389 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_44_401 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_44_41 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_44_413 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_44_419 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_44_421 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_44_433 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_44_445 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_44_457 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_44_469 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_44_475 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_44_477 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_44_489 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_44_501 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_44_513 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_44_53 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_44_65 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_44_77 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_44_83 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_44_85 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_44_97 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_45_105 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_45_111 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_45_113 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_45_125 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_45_137 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_45_149 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_45_15 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_45_161 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_45_167 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_45_169 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_45_181 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_45_193 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_45_205 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_45_217 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_45_223 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_45_225 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_45_237 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_45_249 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_45_261 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_45_27 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_45_273 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_45_279 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_45_281 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_45_293 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_45_3 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_45_305 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_45_317 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_45_329 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_45_335 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_45_337 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_45_349 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_45_361 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_45_373 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_45_385 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_45_39 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_45_391 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_45_393 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_45_405 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_45_417 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_45_429 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_45_441 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_45_447 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_45_449 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_45_461 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_45_473 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_45_485 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_45_497 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_45_503 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_8 FILLER_45_505 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_4 FILLER_45_51 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_45_513 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_45_55 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_45_57 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_45_69 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_45_81 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_45_93 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_46_109 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_46_121 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_46_133 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_46_139 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_46_141 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_46_15 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_46_153 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_46_165 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_46_177 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_46_189 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_46_195 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_46_197 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_46_209 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_46_221 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_46_233 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_46_245 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_46_251 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_46_253 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_46_265 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_46_27 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_46_277 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_46_289 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_46_29 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_46_3 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_46_301 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_46_307 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_46_309 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_46_321 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_46_333 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_46_345 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_46_357 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_46_363 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_46_365 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_46_377 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_46_389 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_46_401 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_46_41 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_46_413 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_46_419 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_46_421 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_46_433 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_46_445 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_46_457 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_46_469 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_46_475 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_46_477 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_46_489 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_46_501 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_46_513 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_46_53 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_46_65 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_46_77 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_46_83 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_46_85 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_46_97 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_47_105 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_47_111 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_47_113 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_47_125 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_47_137 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_47_149 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_47_15 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_47_161 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_47_167 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_47_169 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_47_181 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_47_193 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_47_205 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_47_217 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_47_223 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_47_225 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_47_237 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_47_249 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_47_261 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_47_27 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_47_273 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_47_279 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_47_281 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_47_293 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_47_3 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_47_305 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_47_317 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_47_329 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_47_335 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_47_337 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_47_349 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_47_361 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_47_373 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_47_385 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_47_39 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_47_391 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_47_393 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_47_405 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_47_417 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_47_429 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_47_441 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_47_447 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_47_449 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_47_461 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_47_473 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_47_485 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_47_497 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_47_503 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_8 FILLER_47_505 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_4 FILLER_47_51 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_47_513 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_47_55 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_47_57 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_47_69 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_47_81 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_47_93 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_48_109 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_48_121 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_48_133 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_48_139 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_48_141 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_48_15 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_48_153 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_48_165 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_48_177 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_48_189 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_48_195 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_48_197 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_48_209 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_48_221 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_48_233 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_48_245 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_48_251 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_48_253 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_48_265 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_48_27 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_48_277 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_48_289 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_48_29 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_48_3 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_48_301 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_48_307 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_48_309 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_48_321 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_48_333 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_48_345 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_48_357 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_48_363 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_48_365 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_48_377 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_48_389 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_48_401 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_48_41 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_48_413 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_48_419 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_48_421 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_48_433 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_48_445 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_48_457 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_48_469 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_48_475 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_48_477 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_48_489 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_48_501 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_48_513 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_48_53 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_48_65 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_48_77 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_48_83 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_48_85 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_48_97 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_49_105 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_49_111 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_49_113 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_49_125 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_49_137 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_49_149 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_49_15 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_49_161 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_49_167 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_49_169 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_49_181 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_49_193 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_49_205 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_49_217 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_49_223 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_49_225 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_49_237 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_49_249 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_49_261 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_49_27 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_49_273 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_49_279 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_49_281 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_49_293 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_49_3 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_49_305 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_49_317 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_49_329 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_49_335 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_49_337 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_49_349 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_49_361 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_49_373 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_49_385 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_49_39 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_49_391 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_49_393 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_49_405 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_49_417 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_49_429 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_49_441 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_49_447 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_49_449 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_49_461 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_49_473 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_49_485 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_49_497 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_49_503 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_8 FILLER_49_505 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_4 FILLER_49_51 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_49_513 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_49_55 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_49_57 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_49_69 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_49_81 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_49_93 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_4_109 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_4_121 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_4_133 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_4_139 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_4_141 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_4_15 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_4_153 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_4_165 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_4_177 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_4_189 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_4_195 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_4_197 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_4_209 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_4_221 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_4_233 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_4_245 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_4_251 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_4_253 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_4_265 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_4_27 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_4_277 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_4_289 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_4_29 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_4_3 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_4_301 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_4_307 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_4_309 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_4_321 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_4_333 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_4_345 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_4_357 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_4_363 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_4_365 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_4_377 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_4_389 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_4_401 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_4_41 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_4_413 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_4_419 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_4_421 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_4_433 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_4_445 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_4_457 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_4_469 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_4_475 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_4_477 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_4_489 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_4_501 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_4_513 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_4_53 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_4_65 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_4_77 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_4_83 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_4_85 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_4_97 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_50_109 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_50_121 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_50_133 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_50_139 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_50_141 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_50_15 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_50_153 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_50_165 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_50_177 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_50_189 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_50_195 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_50_197 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_50_209 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_50_221 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_50_233 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_50_245 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_50_251 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_50_253 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_50_265 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_50_27 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_50_277 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_50_289 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_50_29 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_50_3 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_50_301 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_50_307 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_50_309 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_50_321 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_50_333 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_50_345 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_50_357 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_50_363 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_50_365 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_50_377 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_50_389 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_50_401 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_50_41 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_50_413 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_50_419 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_50_421 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_50_433 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_50_445 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_50_457 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_50_469 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_50_475 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_50_477 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_50_489 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_50_501 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_50_513 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_50_53 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_50_65 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_50_77 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_50_83 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_50_85 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_50_97 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_51_105 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_51_111 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_51_113 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_51_125 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_51_137 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_51_149 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_51_15 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_51_161 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_51_167 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_51_169 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_51_181 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_51_193 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_51_205 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_51_217 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_51_223 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_51_225 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_51_237 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_51_249 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_51_261 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_51_27 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_51_273 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_51_279 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_51_281 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_51_293 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_51_3 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_51_305 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_51_317 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_51_329 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_51_335 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_51_337 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_51_349 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_51_361 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_51_373 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_51_385 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_51_39 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_51_391 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_51_393 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_51_405 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_51_417 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_51_429 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_51_441 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_51_447 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_51_449 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_51_461 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_51_473 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_51_485 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_51_497 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_51_503 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_8 FILLER_51_505 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_4 FILLER_51_51 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_51_513 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_51_55 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_51_57 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_51_69 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_51_81 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_51_93 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_52_109 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_52_121 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_52_133 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_52_139 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_52_141 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_52_15 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_52_153 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_52_165 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_52_177 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_52_189 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_52_195 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_52_197 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_52_209 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_52_221 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_52_233 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_52_245 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_52_251 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_52_253 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_52_265 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_52_27 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_52_277 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_52_289 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_52_29 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_52_3 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_52_301 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_52_307 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_52_309 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_52_321 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_52_333 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_52_345 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_52_357 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_52_363 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_52_365 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_52_377 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_52_389 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_52_401 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_52_41 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_52_413 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_52_419 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_52_421 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_52_433 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_52_445 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_52_457 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_52_469 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_52_475 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_52_477 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_52_489 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_52_501 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_52_513 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_52_53 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_52_65 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_52_77 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_52_83 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_52_85 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_52_97 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_53_105 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_53_111 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_53_113 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_53_125 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_53_137 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_53_149 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_53_15 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_53_161 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_53_167 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_53_169 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_53_181 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_53_193 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_53_205 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_53_217 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_53_223 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_53_225 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_53_237 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_53_249 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_53_261 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_53_27 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_53_273 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_53_279 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_53_281 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_53_293 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_53_3 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_53_305 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_53_317 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_53_329 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_53_335 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_53_337 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_53_349 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_53_361 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_53_373 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_53_385 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_53_39 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_53_391 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_53_393 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_53_405 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_53_417 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_53_429 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_53_441 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_53_447 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_53_449 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_53_461 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_53_473 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_53_485 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_53_497 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_53_503 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_8 FILLER_53_505 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_4 FILLER_53_51 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_53_513 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_53_55 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_53_57 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_53_69 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_53_81 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_53_93 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_54_109 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_54_121 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_54_133 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_54_139 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_54_141 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_54_15 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_54_153 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_54_165 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_54_177 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_54_189 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_54_195 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_54_197 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_54_209 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_54_221 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_54_233 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_54_245 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_54_251 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_54_253 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_54_265 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_54_27 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_54_277 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_54_289 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_54_29 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_54_3 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_54_301 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_54_307 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_54_309 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_54_321 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_54_333 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_54_345 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_54_357 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_54_363 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_54_365 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_54_377 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_54_389 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_54_401 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_54_41 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_54_413 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_54_419 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_54_421 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_54_433 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_54_445 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_54_457 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_54_469 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_54_475 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_54_477 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_54_489 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_54_501 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_54_513 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_54_53 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_54_65 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_54_77 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_54_83 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_54_85 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_54_97 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_55_105 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_55_111 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_55_113 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_55_125 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_55_137 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_55_149 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_55_15 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_55_161 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_55_167 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_55_169 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_55_181 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_55_193 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_55_205 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_55_217 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_55_223 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_55_225 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_55_237 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_55_249 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_55_261 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_55_27 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_55_273 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_55_279 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_55_281 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_55_293 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_55_3 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_55_305 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_55_317 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_55_329 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_55_335 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_55_337 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_55_349 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_55_361 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_55_373 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_55_385 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_55_39 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_55_391 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_55_393 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_55_405 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_55_417 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_55_429 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_55_441 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_55_447 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_55_449 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_55_461 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_55_473 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_55_485 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_55_497 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_55_503 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_8 FILLER_55_505 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_4 FILLER_55_51 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_55_513 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_55_55 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_55_57 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_55_69 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_55_81 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_55_93 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_56_109 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_56_121 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_56_133 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_56_139 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_56_141 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_56_15 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_56_153 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_56_165 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_56_177 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_56_189 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_56_195 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_56_197 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_56_209 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_56_221 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_56_233 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_56_245 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_56_251 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_56_253 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_56_265 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_56_27 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_56_277 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_56_289 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_56_29 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_56_3 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_56_301 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_56_307 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_56_309 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_56_321 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_56_333 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_56_345 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_56_357 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_56_363 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_56_365 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_56_377 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_56_389 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_56_401 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_56_41 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_56_413 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_56_419 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_56_421 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_56_433 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_56_445 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_56_457 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_56_469 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_56_475 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_56_477 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_56_489 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_56_501 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_56_513 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_56_53 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_56_65 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_56_77 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_56_83 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_56_85 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_56_97 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_57_105 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_57_111 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_57_113 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_57_125 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_57_137 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_57_149 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_57_15 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_57_161 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_57_167 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_57_169 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_57_181 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_57_193 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_57_205 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_57_217 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_57_223 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_57_225 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_57_237 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_57_249 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_57_261 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_57_27 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_57_273 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_57_279 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_57_281 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_57_293 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_57_3 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_57_305 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_57_317 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_57_329 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_57_335 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_57_337 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_57_349 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_57_361 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_57_373 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_57_385 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_57_39 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_57_391 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_57_393 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_57_405 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_57_417 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_57_429 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_57_441 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_57_447 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_57_449 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_57_461 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_57_473 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_57_485 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_57_497 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_57_503 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_8 FILLER_57_505 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_4 FILLER_57_51 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_57_513 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_57_55 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_57_57 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_57_69 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_57_81 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_57_93 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_58_109 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_58_121 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_58_133 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_58_139 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_58_141 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_58_15 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_58_153 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_58_165 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_58_177 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_58_189 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_58_195 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_58_197 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_58_209 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_58_221 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_58_233 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_58_245 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_58_251 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_58_253 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_58_265 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_58_27 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_58_277 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_58_289 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_58_29 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_58_3 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_58_301 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_58_307 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_58_309 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_58_321 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_58_333 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_58_345 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_58_357 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_58_363 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_58_365 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_58_377 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_58_389 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_58_401 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_58_41 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_58_413 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_58_419 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_58_421 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_58_433 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_58_445 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_58_457 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_58_469 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_58_475 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_58_477 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_58_489 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_58_501 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_58_513 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_58_53 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_58_65 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_58_77 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_58_83 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_58_85 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_58_97 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_59_105 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_59_111 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_59_113 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_59_125 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_59_137 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_59_149 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_59_15 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_59_161 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_59_167 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_59_169 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_59_181 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_59_193 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_59_205 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_59_217 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_59_223 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_59_225 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_59_237 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_59_249 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_59_261 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_59_27 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_59_273 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_59_279 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_59_281 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_59_293 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_59_3 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_59_305 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_59_317 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_59_329 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_59_335 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_59_337 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_59_349 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_59_361 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_59_373 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_59_385 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_59_39 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_59_391 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_59_393 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_59_405 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_59_417 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_59_429 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_59_441 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_59_447 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_59_449 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_59_461 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_59_473 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_59_485 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_59_497 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_59_503 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_8 FILLER_59_505 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_4 FILLER_59_51 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_59_513 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_59_55 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_59_57 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_59_69 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_59_81 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_59_93 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_5_105 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_5_111 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_5_113 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_5_125 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_5_137 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_5_149 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_5_15 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_5_161 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_5_167 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_5_169 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_5_181 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_5_193 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_5_205 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_5_217 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_5_223 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_5_225 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_5_237 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_5_249 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_5_261 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_5_27 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_5_273 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_5_279 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_5_281 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_5_293 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_5_3 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_5_305 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_5_317 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_5_329 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_5_335 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_5_337 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_5_349 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_5_361 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_5_373 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_5_385 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_5_39 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_5_391 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_5_393 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_5_405 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_5_417 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_5_429 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_5_441 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_5_447 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_5_449 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_5_461 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_5_473 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_5_485 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_5_497 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_5_503 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_8 FILLER_5_505 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_4 FILLER_5_51 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_5_513 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_5_55 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_5_57 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_5_69 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_5_81 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_5_93 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_60_109 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_60_121 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_60_133 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_60_139 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_60_141 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_60_15 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_60_153 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_60_165 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_60_177 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_60_189 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_60_195 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_60_197 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_60_209 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_60_221 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_60_233 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_60_245 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_60_251 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_60_253 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_60_265 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_60_27 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_60_277 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_60_289 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_60_29 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_60_3 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_60_301 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_60_307 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_60_309 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_60_321 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_60_333 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_60_345 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_60_357 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_60_363 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_60_365 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_60_377 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_60_389 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_60_401 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_60_41 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_60_413 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_60_419 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_60_421 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_60_433 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_60_445 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_60_457 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_60_469 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_60_475 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_60_477 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_60_489 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_60_501 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_60_513 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_60_53 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_60_65 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_60_77 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_60_83 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_60_85 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_60_97 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_61_105 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_61_111 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_61_113 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_61_125 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_61_137 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_61_149 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_61_15 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_61_161 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_61_167 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_61_169 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_61_181 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_61_193 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_61_205 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_61_217 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_61_223 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_61_225 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_61_237 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_61_249 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_61_261 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_61_27 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_61_273 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_61_279 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_61_281 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_61_293 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_61_3 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_61_305 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_61_317 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_61_329 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_61_335 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_61_337 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_61_349 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_61_361 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_61_373 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_61_385 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_61_39 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_61_391 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_61_393 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_61_405 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_61_417 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_61_429 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_61_441 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_61_447 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_61_449 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_61_461 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_61_473 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_61_485 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_61_497 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_61_503 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_8 FILLER_61_505 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_4 FILLER_61_51 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_61_513 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_61_55 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_61_57 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_61_69 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_61_81 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_61_93 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_62_109 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_62_121 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_62_133 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_62_139 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_62_141 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_62_15 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_62_153 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_62_165 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_62_177 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_62_189 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_62_195 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_62_197 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_62_209 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_62_221 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_62_233 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_62_245 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_62_251 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_62_253 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_62_265 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_62_27 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_62_277 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_62_289 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_62_29 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_62_3 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_62_301 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_62_307 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_62_309 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_62_321 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_62_333 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_62_345 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_62_357 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_62_363 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_62_365 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_62_377 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_62_389 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_62_401 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_62_41 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_62_413 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_62_419 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_62_421 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_62_433 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_62_445 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_62_457 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_62_469 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_62_475 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_62_477 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_62_489 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_62_501 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_62_513 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_62_53 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_62_65 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_62_77 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_62_83 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_62_85 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_62_97 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_63_105 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_63_111 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_63_113 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_63_125 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_63_137 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_63_149 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_63_15 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_63_161 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_63_167 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_63_169 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_63_181 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_63_193 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_63_205 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_63_217 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_63_223 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_63_225 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_63_237 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_63_249 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_63_261 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_63_27 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_63_273 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_63_279 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_63_281 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_63_293 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_63_3 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_63_305 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_63_317 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_63_329 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_63_335 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_63_337 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_63_349 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_63_361 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_63_373 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_63_385 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_63_39 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_63_391 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_63_393 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_63_405 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_63_417 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_63_429 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_63_441 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_63_447 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_63_449 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_63_461 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_63_473 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_63_485 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_63_497 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_63_503 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_8 FILLER_63_505 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_4 FILLER_63_51 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_63_513 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_63_55 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_63_57 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_63_69 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_63_81 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_63_93 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_64_109 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_64_121 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_64_133 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_64_139 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_64_141 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_64_15 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_64_153 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_64_165 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_64_177 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_64_189 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_64_195 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_64_197 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_64_209 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_64_221 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_64_233 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_64_245 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_64_251 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_64_253 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_64_265 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_64_27 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_64_277 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_64_289 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_64_29 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_64_3 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_64_301 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_64_307 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_64_309 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_64_321 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_64_333 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_64_345 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_64_357 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_64_363 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_64_365 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_64_377 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_64_389 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_64_401 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_64_41 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_64_413 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_64_419 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_64_421 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_64_433 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_64_445 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_64_457 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_64_469 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_64_475 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_64_477 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_64_489 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_64_501 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_64_513 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_64_53 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_64_65 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_64_77 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_64_83 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_64_85 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_64_97 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_65_105 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_65_111 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_65_113 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_65_125 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_65_137 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_65_149 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_65_15 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_65_161 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_65_167 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_65_169 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_65_181 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_65_193 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_65_205 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_65_217 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_65_223 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_65_225 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_65_237 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_65_249 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_65_261 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_65_27 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_65_273 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_65_279 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_65_281 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_65_293 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_65_3 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_65_305 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_65_317 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_65_329 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_65_335 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_65_337 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_65_349 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_65_361 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_65_373 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_65_385 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_65_39 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_65_391 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_65_393 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_65_405 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_65_417 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_65_429 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_65_441 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_65_447 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_65_449 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_65_461 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_65_473 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_65_485 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_65_497 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_65_503 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_8 FILLER_65_505 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_4 FILLER_65_51 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_65_513 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_65_55 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_65_57 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_65_69 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_65_81 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_65_93 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_66_109 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_66_121 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_66_133 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_66_139 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_66_141 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_66_15 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_66_153 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_66_165 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_66_177 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_66_189 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_66_195 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_66_197 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_66_209 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_66_221 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_66_233 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_66_245 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_66_251 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_66_253 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_66_265 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_66_27 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_66_277 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_66_289 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_66_29 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_66_3 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_66_301 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_66_307 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_66_309 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_66_321 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_66_333 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_66_345 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_66_357 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_66_363 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_66_365 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_66_377 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_66_389 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_66_401 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_66_41 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_66_413 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_66_419 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_66_421 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_66_433 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_66_445 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_66_457 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_66_469 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_66_475 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_66_477 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_66_489 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_66_501 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_66_513 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_66_53 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_66_65 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_66_77 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_66_83 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_66_85 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_66_97 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_67_105 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_67_111 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_67_113 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_67_125 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_67_137 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_67_149 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_67_15 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_67_161 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_67_167 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_67_169 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_67_181 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_67_193 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_67_205 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_67_217 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_67_223 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_67_225 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_67_237 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_67_249 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_67_261 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_67_27 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_67_273 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_67_279 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_67_281 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_67_293 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_67_3 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_67_305 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_67_317 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_67_329 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_67_335 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_67_337 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_67_349 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_67_361 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_67_373 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_67_385 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_67_39 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_67_391 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_67_393 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_67_405 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_67_417 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_67_429 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_67_441 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_67_447 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_67_449 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_67_461 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_67_473 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_67_485 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_67_497 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_67_503 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_8 FILLER_67_505 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_4 FILLER_67_51 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_67_513 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_67_55 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_67_57 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_67_69 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_67_81 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_67_93 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_68_109 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_68_121 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_68_133 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_68_139 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_68_141 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_68_15 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_68_153 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_68_165 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_68_177 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_68_189 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_68_195 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_68_197 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_68_209 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_68_221 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_68_233 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_68_245 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_68_251 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_68_253 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_68_265 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_68_27 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_68_277 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_68_289 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_68_29 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_68_3 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_68_301 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_68_307 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_68_309 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_68_321 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_68_333 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_68_345 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_68_357 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_68_363 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_68_365 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_68_377 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_68_389 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_68_401 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_68_41 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_68_413 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_68_419 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_68_421 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_68_433 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_68_445 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_68_457 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_68_469 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_68_475 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_68_477 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_68_489 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_68_501 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_68_513 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_68_53 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_68_65 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_68_77 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_68_83 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_68_85 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_68_97 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_69_105 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_69_111 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_69_113 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_69_125 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_69_137 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_69_149 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_69_15 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_69_161 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_69_167 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_69_169 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_69_181 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_69_193 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_69_205 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_69_217 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_69_223 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_69_225 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_69_237 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_69_249 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_69_261 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_69_27 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_69_273 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_69_279 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_69_281 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_69_293 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_69_3 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_69_305 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_69_317 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_69_329 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_69_335 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_69_337 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_69_349 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_69_361 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_69_373 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_69_385 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_69_39 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_69_391 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_69_393 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_69_405 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_69_417 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_69_429 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_69_441 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_69_447 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_69_449 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_69_461 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_69_473 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_69_485 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_69_497 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_69_503 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_8 FILLER_69_505 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_4 FILLER_69_51 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_69_513 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_69_55 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_69_57 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_69_69 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_69_81 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_69_93 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_6_109 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_6_121 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_6_133 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_6_139 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_6_141 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_6_15 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_6_153 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_6_165 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_6_177 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_6_189 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_6_195 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_6_197 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_6_209 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_6_221 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_6_233 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_6_245 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_6_251 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_6_253 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_6_265 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_6_27 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_6_277 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_6_289 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_6_29 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_6_3 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_6_301 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_6_307 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_6_309 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_6_321 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_6_333 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_6_345 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_6_357 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_6_363 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_6_365 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_6_377 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_6_389 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_6_401 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_6_41 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_6_413 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_6_419 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_6_421 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_6_433 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_6_445 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_6_457 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_6_469 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_6_475 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_6_477 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_6_489 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_6_501 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_6_513 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_6_53 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_6_65 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_6_77 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_6_83 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_6_85 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_6_97 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_70_109 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_70_121 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_70_133 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_70_139 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_70_141 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_70_15 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_70_153 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_70_165 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_70_177 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_70_189 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_70_195 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_70_197 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_70_209 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_70_221 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_70_233 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_70_245 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_70_251 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_70_253 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_70_265 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_70_27 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_70_277 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_70_289 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_70_29 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_70_3 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_70_301 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_70_307 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_70_309 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_70_321 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_70_333 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_70_345 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_70_357 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_70_363 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_70_365 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_70_377 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_70_389 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_70_401 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_70_41 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_70_413 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_70_419 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_70_421 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_70_433 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_70_445 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_70_457 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_70_469 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_70_475 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_70_477 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_70_489 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_70_501 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_70_513 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_70_53 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_70_65 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_70_77 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_70_83 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_70_85 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_70_97 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_71_105 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_71_111 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_71_113 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_71_125 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_71_137 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_71_149 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_71_15 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_71_161 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_71_167 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_71_169 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_71_181 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_71_193 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_71_205 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_71_217 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_71_223 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_71_225 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_71_237 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_71_249 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_71_261 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_71_27 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_71_273 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_71_279 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_71_281 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_71_293 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_71_3 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_71_305 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_71_317 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_71_329 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_71_335 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_71_337 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_71_349 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_71_361 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_71_373 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_71_385 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_71_39 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_71_391 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_71_393 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_71_405 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_71_417 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_71_429 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_71_441 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_71_447 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_71_449 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_71_461 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_71_473 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_71_485 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_71_497 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_71_503 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_8 FILLER_71_505 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_4 FILLER_71_51 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_71_513 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_71_55 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_71_57 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_71_69 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_71_81 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_71_93 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_72_109 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_72_121 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_72_133 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_72_139 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_72_141 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_72_15 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_72_153 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_72_165 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_72_177 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_72_189 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_72_195 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_72_197 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_72_209 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_72_221 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_72_233 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_72_245 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_72_251 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_72_253 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_72_265 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_72_27 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_72_277 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_72_289 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_72_29 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_72_3 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_72_301 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_72_307 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_72_309 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_72_321 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_72_333 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_72_345 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_72_357 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_72_363 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_72_365 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_72_377 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_72_389 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_72_401 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_72_41 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_72_413 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_72_419 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_72_421 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_72_433 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_72_445 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_72_457 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_72_469 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_72_475 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_72_477 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_72_489 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_72_501 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_72_513 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_72_53 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_72_65 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_72_77 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_72_83 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_72_85 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_72_97 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_73_105 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_73_111 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_73_113 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_73_125 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_73_137 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_73_149 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_73_15 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_73_161 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_73_167 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_73_169 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_73_181 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_73_193 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_73_205 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_73_217 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_73_223 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_73_225 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_73_237 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_73_249 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_73_261 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_73_27 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_73_273 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_73_279 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_73_281 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_73_293 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_73_3 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_73_305 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_73_317 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_73_329 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_73_335 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_73_337 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_73_349 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_73_361 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_73_373 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_73_385 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_73_39 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_73_391 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_73_393 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_73_405 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_73_417 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_73_429 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_73_441 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_73_447 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_73_449 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_73_461 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_73_473 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_73_485 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_73_497 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_73_503 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_8 FILLER_73_505 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_4 FILLER_73_51 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_73_513 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_73_55 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_73_57 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_73_69 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_73_81 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_73_93 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_74_109 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_74_121 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_74_133 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_74_139 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_74_141 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_74_15 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_74_153 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_74_165 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_74_177 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_74_189 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_74_195 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_74_197 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_74_209 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_74_221 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_74_233 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_74_245 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_74_251 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_74_253 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_74_265 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_74_27 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_74_277 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_74_289 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_74_29 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_74_3 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_74_301 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_74_307 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_74_309 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_74_321 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_74_333 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_74_345 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_74_357 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_74_363 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_74_365 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_74_377 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_74_389 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_74_401 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_74_41 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_74_413 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_74_419 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_74_421 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_74_433 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_74_445 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_74_457 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_74_469 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_74_475 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_74_477 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_74_489 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_74_501 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_74_513 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_74_53 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_74_65 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_74_77 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_74_83 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_74_85 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_74_97 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_75_105 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_75_111 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_75_113 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_75_125 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_75_137 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_75_149 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_75_15 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_75_161 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_75_167 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_75_169 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_75_181 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_75_193 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_75_205 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_75_217 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_75_223 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_75_225 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_75_237 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_75_249 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_75_261 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_75_27 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_75_273 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_75_279 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_75_281 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_75_293 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_75_3 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_75_305 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_75_317 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_75_329 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_75_335 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_75_337 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_75_349 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_75_361 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_75_373 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_75_385 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_75_39 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_75_391 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_75_393 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_75_405 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_75_417 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_75_429 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_75_441 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_75_447 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_75_449 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_75_461 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_75_473 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_75_485 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_75_497 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_75_503 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_8 FILLER_75_505 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_4 FILLER_75_51 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_75_513 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_75_55 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_75_57 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_75_69 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_75_81 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_75_93 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_76_109 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_76_121 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_76_133 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_76_139 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_76_141 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_76_15 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_76_153 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_76_165 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_76_177 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_76_189 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_76_195 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_76_197 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_76_209 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_76_221 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_76_233 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_76_245 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_76_251 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_76_253 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_76_265 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_76_27 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_76_277 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_76_289 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_76_29 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_76_3 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_76_301 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_76_307 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_76_309 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_76_321 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_76_333 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_76_345 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_76_357 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_76_363 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_76_365 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_76_377 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_76_389 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_76_401 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_76_41 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_76_413 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_76_419 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_76_421 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_76_433 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_76_445 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_76_457 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_76_469 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_76_475 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_76_477 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_76_489 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_76_501 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_76_513 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_76_53 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_76_65 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_76_77 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_76_83 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_76_85 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_76_97 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_77_105 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_77_111 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_77_113 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_77_125 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_77_137 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_77_149 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_77_15 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_77_161 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_77_167 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_77_169 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_77_181 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_77_193 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_77_205 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_77_217 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_77_223 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_77_225 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_77_237 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_77_249 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_77_261 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_77_27 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_77_273 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_77_279 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_77_281 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_77_293 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_77_3 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_77_305 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_77_317 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_77_329 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_77_335 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_77_337 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_77_349 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_77_361 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_77_373 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_77_385 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_77_39 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_77_391 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_77_393 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_77_405 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_77_417 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_77_429 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_77_441 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_77_447 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_77_449 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_77_461 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_77_473 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_77_485 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_77_497 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_77_503 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_8 FILLER_77_505 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_4 FILLER_77_51 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_77_513 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_77_55 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_77_57 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_77_69 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_77_81 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_77_93 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_78_109 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_78_121 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_78_133 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_78_139 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_78_141 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_78_15 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_78_153 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_78_165 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_78_177 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_78_189 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_78_195 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_78_197 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_78_209 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_78_221 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_78_233 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_78_245 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_78_251 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_78_253 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_78_265 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_78_27 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_78_277 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_78_289 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_78_29 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_78_3 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_78_301 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_78_307 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_78_309 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_78_321 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_78_333 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_78_345 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_78_357 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_78_363 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_78_365 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_78_377 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_78_389 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_78_401 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_78_41 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_78_413 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_78_419 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_78_421 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_78_433 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_78_445 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_78_457 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_78_469 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_78_475 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_78_477 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_78_489 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_78_501 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_78_513 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_78_53 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_78_65 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_78_77 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_78_83 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_78_85 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_78_97 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_79_105 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_79_111 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_79_113 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_79_125 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_79_137 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_79_149 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_79_15 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_79_161 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_79_167 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_79_169 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_79_181 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_79_193 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_79_205 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_79_217 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_79_223 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_79_225 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_79_237 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_79_249 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_79_261 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_79_27 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_79_273 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_79_279 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_79_281 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_79_293 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_79_3 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_79_305 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_79_317 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_79_329 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_79_335 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_79_337 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_79_349 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_79_361 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_79_373 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_79_385 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_79_39 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_79_391 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_79_393 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_79_405 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_79_417 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_79_429 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_79_441 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_79_447 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_79_449 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_79_461 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_79_473 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_79_485 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_79_497 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_79_503 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_8 FILLER_79_505 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_4 FILLER_79_51 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_79_513 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_79_55 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_79_57 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_79_69 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_79_81 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_79_93 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_7_105 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_7_111 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_7_113 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_7_125 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_7_137 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_7_149 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_7_15 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_7_161 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_7_167 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_7_169 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_7_181 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_7_193 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_7_205 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_7_217 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_7_223 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_7_225 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_7_237 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_7_249 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_7_261 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_7_27 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_7_273 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_7_279 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_7_281 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_7_293 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_7_3 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_7_305 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_7_317 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_7_329 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_7_335 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_7_337 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_7_349 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_7_361 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_7_373 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_7_385 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_7_39 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_7_391 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_7_393 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_7_405 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_7_417 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_7_429 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_7_441 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_7_447 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_7_449 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_7_461 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_7_473 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_7_485 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_7_497 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_7_503 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_8 FILLER_7_505 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_4 FILLER_7_51 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_7_513 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_7_55 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_7_57 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_7_69 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_7_81 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_7_93 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_80_109 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_80_121 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_80_133 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_80_139 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_80_141 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_80_15 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_80_153 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_80_165 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_80_177 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_80_189 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_80_195 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_80_197 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_80_209 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_80_221 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_80_233 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_80_245 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_80_251 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_80_253 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_80_265 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_80_27 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_80_277 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_80_289 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_80_29 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_80_3 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_80_301 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_80_307 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_80_309 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_80_321 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_80_333 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_80_345 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_80_357 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_80_363 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_80_365 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_80_377 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_80_389 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_80_401 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_80_41 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_80_413 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_80_419 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_80_421 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_80_433 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_80_445 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_80_457 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_80_469 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_80_475 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_80_477 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_80_489 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_80_501 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_80_513 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_80_53 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_80_65 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_80_77 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_80_83 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_80_85 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_80_97 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_81_105 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_81_111 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_81_113 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_81_125 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_81_137 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_81_149 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_81_15 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_81_161 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_81_167 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_81_169 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_81_181 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_81_193 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_81_205 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_81_217 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_81_223 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_81_225 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_81_237 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_81_249 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_81_261 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_81_27 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_81_273 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_81_279 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_81_281 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_81_293 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_81_3 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_81_305 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_81_317 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_81_329 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_81_335 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_81_337 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_81_349 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_81_361 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_81_373 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_81_385 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_81_39 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_81_391 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_81_393 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_81_405 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_81_417 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_81_429 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_81_441 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_81_447 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_81_449 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_81_461 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_81_473 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_81_485 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_81_497 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_81_503 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_8 FILLER_81_505 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_4 FILLER_81_51 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_81_513 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_81_55 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_81_57 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_81_69 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_81_81 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_81_93 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_82_109 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_82_121 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_82_133 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_82_139 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_82_141 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_82_15 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_82_153 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_82_165 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_82_177 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_82_189 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_82_195 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_82_197 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_82_209 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_82_221 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_82_233 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_82_245 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_82_251 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_82_253 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_82_265 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_82_27 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_82_277 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_82_289 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_82_29 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_82_3 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_82_301 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_82_307 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_82_309 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_82_321 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_82_333 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_82_345 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_82_357 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_82_363 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_82_365 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_82_377 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_82_389 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_82_401 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_82_41 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_82_413 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_82_419 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_82_421 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_82_433 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_82_445 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_82_457 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_82_469 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_82_475 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_82_477 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_82_489 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_82_501 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_82_513 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_82_53 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_82_65 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_82_77 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_82_83 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_82_85 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_82_97 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_83_105 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_83_111 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_83_113 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_83_125 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_83_137 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_83_149 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_83_15 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_83_161 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_83_167 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_83_169 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_83_181 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_83_193 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_83_205 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_83_217 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_83_223 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_83_225 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_83_237 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_83_249 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_83_261 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_83_27 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_83_273 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_83_279 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_83_281 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_83_293 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_83_3 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_83_305 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_83_317 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_83_329 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_83_335 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_83_337 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_83_349 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_83_361 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_83_373 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_83_385 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_83_39 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_83_391 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_83_393 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_83_405 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_83_417 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_83_429 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_83_441 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_83_447 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_83_449 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_83_461 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_83_473 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_83_485 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_83_497 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_83_503 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_8 FILLER_83_505 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_4 FILLER_83_51 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_83_513 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_83_55 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_83_57 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_83_69 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_83_81 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_83_93 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_84_109 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_84_121 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_84_133 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_84_139 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_84_141 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_84_15 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_84_153 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_84_165 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_84_177 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_84_189 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_84_195 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_84_197 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_84_209 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_84_221 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_84_233 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_84_245 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_84_251 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_84_253 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_84_265 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_84_27 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_84_277 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_84_289 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_84_29 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_84_3 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_84_301 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_84_307 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_84_309 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_84_321 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_84_333 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_84_345 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_84_357 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_84_363 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_84_365 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_84_377 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_84_389 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_84_401 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_84_41 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_84_413 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_84_419 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_84_421 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_84_433 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_84_445 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_84_457 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_84_469 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_84_475 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_84_477 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_84_489 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_84_501 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_84_513 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_84_53 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_84_65 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_84_77 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_84_83 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_84_85 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_84_97 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_85_105 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_85_111 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_85_113 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_85_125 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_85_137 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_85_149 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_85_15 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_85_161 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_85_167 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_85_169 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_85_181 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_85_193 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_85_205 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_85_217 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_85_223 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_85_225 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_85_237 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_85_249 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_85_261 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_85_27 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_85_273 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_85_279 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_85_281 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_85_293 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_85_3 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_85_305 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_85_317 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_85_329 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_85_335 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_85_337 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_85_349 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_85_361 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_85_373 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_85_385 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_85_39 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_85_391 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_85_393 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_85_405 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_85_417 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_85_429 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_85_441 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_85_447 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_85_449 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_85_461 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_85_473 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_85_485 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_85_497 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_85_503 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_8 FILLER_85_505 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_4 FILLER_85_51 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_85_513 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_85_55 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_85_57 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_85_69 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_85_81 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_85_93 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_86_109 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_86_121 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_86_133 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_86_139 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_86_141 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_86_15 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_86_153 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_86_165 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_86_177 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_86_189 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_86_195 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_86_197 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_86_209 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_86_221 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_86_233 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_86_245 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_86_251 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_86_253 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_86_265 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_86_27 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_86_277 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_86_289 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_86_29 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_86_3 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_86_301 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_86_307 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_86_309 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_86_321 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_86_333 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_86_345 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_86_357 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_86_363 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_86_365 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_86_377 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_86_389 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_86_401 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_86_41 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_86_413 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_86_419 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_86_421 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_86_433 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_86_445 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_86_457 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_86_469 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_86_475 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_86_477 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_86_489 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_86_501 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_86_513 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_86_53 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_86_65 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_86_77 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_86_83 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_86_85 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_86_97 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_87_105 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_87_111 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_87_113 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_87_125 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_87_137 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_87_149 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_87_15 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_87_161 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_87_167 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_87_169 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_87_181 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_87_193 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_87_205 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_87_217 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_87_223 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_87_225 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_87_237 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_87_249 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_87_261 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_87_27 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_87_273 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_87_279 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_87_281 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_87_293 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_87_3 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_87_305 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_87_317 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_87_329 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_87_335 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_87_337 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_87_349 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_87_361 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_87_373 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_87_385 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_87_39 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_87_391 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_87_393 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_87_405 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_87_417 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_87_429 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_87_441 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_87_447 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_87_449 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_87_461 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_87_473 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_87_485 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_87_497 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_87_503 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_8 FILLER_87_505 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_4 FILLER_87_51 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_87_513 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_87_55 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_87_57 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_87_69 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_87_81 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_87_93 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_88_109 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_88_121 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_88_133 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_88_139 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_88_141 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_88_15 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_88_153 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_88_165 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_88_177 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_88_189 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_88_195 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_88_197 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_88_209 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_88_221 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_88_233 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_88_245 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_88_251 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_88_253 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_88_265 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_88_27 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_88_277 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_88_289 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_88_29 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_88_3 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_88_301 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_88_307 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_88_309 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_88_321 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_88_333 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_88_345 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_88_357 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_88_363 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_88_365 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_88_377 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_88_389 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_88_401 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_88_41 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_88_413 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_88_419 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_88_421 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_88_433 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_88_445 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_88_457 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_88_469 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_88_475 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_88_477 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_88_489 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_88_501 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_88_513 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_88_53 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_88_65 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_88_77 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_88_83 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_88_85 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_88_97 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_89_105 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_89_111 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_89_113 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_89_125 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_89_137 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_89_149 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_89_15 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_89_161 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_89_167 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_89_169 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_89_181 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_89_193 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_89_205 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_89_217 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_89_223 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_89_225 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_89_237 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_89_249 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_89_261 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_89_27 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_89_273 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_89_279 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_89_281 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_89_293 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_89_3 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_89_305 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_89_317 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_89_329 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_89_335 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_89_337 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_89_349 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_89_361 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_89_373 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_89_385 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_89_39 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_89_391 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_89_393 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_89_405 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_89_417 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_89_429 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_89_441 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_89_447 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_89_449 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_89_461 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_89_473 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_89_485 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_89_497 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_89_503 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_8 FILLER_89_505 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_4 FILLER_89_51 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_89_513 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_89_55 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_89_57 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_89_69 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_89_81 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_89_93 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_8_109 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_8_121 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_8_133 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_8_139 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_8_141 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_8_15 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_8_153 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_8_165 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_8_177 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_8_189 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_8_195 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_8_197 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_8_209 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_8_221 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_8_233 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_8_245 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_8_251 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_8_253 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_8_265 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_8_27 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_8_277 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_8_289 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_8_29 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_8_3 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_8_301 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_8_307 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_8_309 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_8_321 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_8_333 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_8_345 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_8_357 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_8_363 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_8_365 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_8_377 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_8_389 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_8_401 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_8_41 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_8_413 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_8_419 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_8_421 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_8_433 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_8_445 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_8_457 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_8_469 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_8_475 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_8_477 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_8_489 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_8_501 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_8_513 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_8_53 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_8_65 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_8_77 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_8_83 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_8_85 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_8_97 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_90_109 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_90_121 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_90_133 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_90_139 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_90_141 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_90_15 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_90_153 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_90_165 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_90_177 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_90_189 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_90_195 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_90_197 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_90_209 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_90_221 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_90_233 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_90_245 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_90_251 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_90_253 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_90_265 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_90_27 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_90_277 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_90_289 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_90_29 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_90_3 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_90_301 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_90_307 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_90_309 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_90_321 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_90_333 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_90_345 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_90_357 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_90_363 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_90_365 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_90_377 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_90_389 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_90_401 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_90_41 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_90_413 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_90_419 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_90_421 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_90_433 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_90_445 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_90_457 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_90_469 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_90_475 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_90_477 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_90_489 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_90_501 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_90_513 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_90_53 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_90_65 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_90_77 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_90_83 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_90_85 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_90_97 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_91_105 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_91_111 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_91_113 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_91_125 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_91_137 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_91_149 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_91_15 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_91_161 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_91_167 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_91_169 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_91_181 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_91_193 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_91_205 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_91_217 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_91_223 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_91_225 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_91_237 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_91_249 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_91_261 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_91_27 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_91_273 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_91_279 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_91_281 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_91_293 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_91_3 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_91_305 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_91_317 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_91_329 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_91_335 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_91_337 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_91_349 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_91_361 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_91_373 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_91_385 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_91_39 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_91_391 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_91_393 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_91_405 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_91_417 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_91_429 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_91_441 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_91_447 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_91_449 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_91_461 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_91_473 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_91_485 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_91_497 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_91_503 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_8 FILLER_91_505 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_4 FILLER_91_51 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_91_513 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_91_55 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_91_57 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_91_69 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_91_81 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_91_93 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_92_109 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_92_121 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_92_133 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_92_139 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_92_141 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_92_15 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_92_153 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_92_165 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_92_177 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_92_189 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_92_195 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_92_197 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_92_209 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_92_221 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_92_233 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_92_245 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_92_251 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_92_253 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_92_265 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_92_27 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_92_277 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_92_289 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_92_29 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_92_3 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_92_301 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_92_307 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_92_309 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_92_321 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_92_333 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_92_345 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_92_357 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_92_363 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_92_365 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_92_377 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_92_389 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_92_401 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_92_41 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_92_413 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_92_419 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_92_421 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_92_433 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_92_445 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_92_457 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_92_469 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_92_475 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_92_477 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_92_489 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_92_501 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_92_513 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_92_53 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_92_65 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_92_77 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_92_83 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_92_85 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_92_97 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_93_105 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_93_111 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_93_113 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_93_125 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_93_137 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_93_149 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_93_15 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_93_161 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_93_167 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_93_169 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_93_181 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_93_193 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_93_205 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_93_217 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_93_223 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_93_225 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_93_237 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_93_249 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_93_261 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_93_27 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_93_273 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_93_279 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_93_281 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_93_293 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_93_3 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_93_305 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_93_317 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_93_329 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_93_335 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_93_337 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_93_349 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_93_361 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_93_373 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_93_385 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_93_39 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_93_391 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_93_393 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_93_405 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_93_417 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_93_429 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_93_441 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_93_447 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_93_449 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_93_461 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_93_473 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_93_485 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_93_497 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_93_503 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_8 FILLER_93_505 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_4 FILLER_93_51 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_93_513 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_93_55 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_93_57 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_93_69 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_93_81 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_93_93 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_94_109 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_94_121 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_94_133 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_94_139 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_94_141 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_94_15 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_94_153 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_94_165 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_94_177 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_94_189 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_94_195 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_94_197 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_94_209 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_94_221 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_94_233 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_94_245 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_94_251 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_94_253 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_94_265 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_94_27 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_94_277 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_94_289 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_94_29 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_94_3 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_94_301 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_94_307 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_94_309 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_94_321 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_94_333 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_94_345 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_94_357 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_94_363 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_94_365 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_94_377 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_94_389 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_94_401 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_94_41 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_94_413 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_94_419 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_94_421 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_94_433 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_94_445 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_94_457 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_94_469 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_94_475 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_94_477 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_94_489 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_94_501 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_94_513 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_94_53 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_94_65 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_94_77 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_94_83 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_94_85 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_94_97 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_95_105 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_95_111 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_95_113 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_95_125 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_95_137 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_95_149 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_95_15 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_95_161 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_95_167 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_95_169 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_95_181 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_95_193 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_95_205 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_95_217 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_95_223 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_95_225 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_95_237 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_95_249 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_95_261 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_95_27 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_95_273 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_95_279 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_95_281 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_95_293 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_95_3 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_95_305 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_95_317 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_95_329 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_95_335 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_95_337 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_95_349 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_95_361 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_95_373 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_95_385 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_95_39 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_95_391 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_95_393 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_95_405 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_95_417 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_95_429 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_95_441 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_95_447 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_95_449 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_95_461 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_95_473 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_95_485 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_95_497 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_95_503 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_8 FILLER_95_505 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_4 FILLER_95_51 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_95_513 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_95_55 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_95_57 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_95_69 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_95_81 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_95_93 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_96_109 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_96_121 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_96_133 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_96_139 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_96_141 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_96_15 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_96_153 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_96_165 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_96_177 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_96_189 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_96_195 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_96_197 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_96_209 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_96_221 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_96_233 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_96_245 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_96_251 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_96_253 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_96_265 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_96_27 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_96_277 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_96_289 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_96_29 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_96_3 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_96_301 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_96_307 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_96_309 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_96_321 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_96_333 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_96_345 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_96_357 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_96_363 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_96_365 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_96_377 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_96_389 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_96_401 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_96_41 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_96_413 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_96_419 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_96_421 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_96_433 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_96_445 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_96_457 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_96_469 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_96_475 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_96_477 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_96_489 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_96_501 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_96_513 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_96_53 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_96_65 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_96_77 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_96_83 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_96_85 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_96_97 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_97_105 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_97_111 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_97_113 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_97_125 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_97_137 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_97_149 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_97_15 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_97_161 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_97_167 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_97_169 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_97_181 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_97_193 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_97_205 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_97_217 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_97_223 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_97_225 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_97_237 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_97_249 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_97_261 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_97_27 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_97_273 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_97_279 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_97_281 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_97_293 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_97_3 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_97_305 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_97_317 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_97_329 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_97_335 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_97_337 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_97_349 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_97_361 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_97_373 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_97_385 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_97_39 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_97_391 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_97_393 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_97_405 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_97_417 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_97_429 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_97_441 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_97_447 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_97_449 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_97_461 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_97_473 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_97_485 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_97_497 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_97_503 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_8 FILLER_97_505 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_4 FILLER_97_51 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_97_513 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_97_55 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_97_57 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_97_69 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_97_81 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_97_93 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_98_109 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_98_121 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_98_133 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_98_139 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_98_141 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_98_15 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_98_153 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_98_165 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_98_177 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_98_189 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_98_195 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_98_197 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_98_209 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_98_221 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_98_233 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_98_245 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_98_251 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_98_253 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_98_265 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_98_27 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_98_277 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_98_289 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_98_29 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_98_3 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_98_301 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_98_307 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_98_309 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_98_321 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_98_333 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_98_345 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_98_357 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_98_363 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_98_365 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_98_377 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_98_389 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_98_401 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_98_41 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_98_413 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_98_419 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_98_421 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_98_433 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_98_445 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_98_457 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_98_469 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_98_475 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_98_477 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_98_489 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_98_501 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_98_513 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_98_53 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_98_65 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_98_77 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_98_83 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_98_85 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_98_97 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_99_105 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_99_111 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_99_113 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_99_125 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_99_137 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_99_149 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_99_15 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_99_161 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_99_167 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_99_169 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_99_181 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_99_193 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_99_205 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_99_217 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_99_223 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_99_225 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_99_237 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_99_249 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_99_261 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_99_27 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_99_273 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_99_279 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_99_281 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_99_293 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_99_3 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_99_305 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_99_317 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_99_329 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_99_335 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_99_337 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_99_349 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_99_361 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_99_373 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_99_385 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_99_39 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_99_391 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_99_393 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_99_405 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_99_417 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_99_429 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_99_441 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_99_447 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_99_449 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_99_461 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_99_473 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_99_485 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_99_497 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_99_503 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_8 FILLER_99_505 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_4 FILLER_99_51 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_99_513 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_99_55 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_99_57 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_99_69 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_99_81 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_99_93 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_9_105 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_9_111 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_9_113 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_9_125 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_9_137 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_9_149 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_9_15 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_9_161 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_9_167 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_9_169 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_9_181 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_9_193 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_9_205 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_9_217 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_9_223 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_9_225 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_9_237 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_9_249 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_9_261 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_9_27 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_9_273 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_9_279 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_9_281 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_9_293 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_9_3 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_9_305 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_9_317 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_9_329 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_9_335 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_9_337 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_9_349 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_9_361 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_9_373 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_9_385 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_9_39 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_9_391 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_9_393 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_9_405 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_9_417 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_9_429 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_9_441 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_9_447 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_9_449 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_9_461 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_9_473 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_9_485 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_6 FILLER_9_497 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_9_503 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_8 FILLER_9_505 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_4 FILLER_9_51 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 FILLER_9_513 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__fill_1 FILLER_9_55 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_9_57 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_9_69 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_9_81 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_ef_sc_hd__decap_12 FILLER_9_93 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_0 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_1 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_10 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_100 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_101 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_102 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_103 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_104 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_105 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_106 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_107 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_108 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_109 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_11 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_110 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_111 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_112 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_113 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_114 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_115 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_116 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_117 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_118 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_119 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_12 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_120 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_121 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_122 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_123 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_124 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_125 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_126 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_127 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_128 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_129 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_13 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_130 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_131 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_132 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_133 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_134 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_135 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_136 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_137 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_138 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_139 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_14 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_140 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_141 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_142 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_143 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_144 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_145 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_146 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_147 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_148 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_149 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_15 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_150 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_151 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_152 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_153 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_154 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_155 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_156 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_157 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_158 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_159 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_16 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_160 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_161 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_162 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_163 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_164 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_165 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_166 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_167 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_168 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_169 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_17 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_170 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_171 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_172 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_173 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_174 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_175 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_176 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_177 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_178 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_179 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_18 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_180 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_181 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_182 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_183 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_184 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_185 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_186 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_187 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_188 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_189 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_19 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_190 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_191 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_192 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_193 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_194 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_195 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_196 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_197 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_198 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_199 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_2 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_20 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_200 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_201 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_202 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_203 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_204 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_205 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_206 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_207 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_208 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_209 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_21 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_210 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_211 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_212 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_213 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_214 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_215 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_216 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_217 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_218 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_219 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_22 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_220 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_221 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_222 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_223 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_224 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_225 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_226 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_227 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_228 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_229 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_23 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_230 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_231 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_232 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_233 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_234 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_235 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_236 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_237 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_238 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_239 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_24 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_240 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_241 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_242 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_243 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_244 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_245 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_246 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_247 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_248 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_249 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_25 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_250 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_251 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_252 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_253 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_254 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_255 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_256 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_257 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_258 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_259 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_26 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_260 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_261 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_262 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_263 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_264 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_265 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_266 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_267 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_268 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_269 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_27 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_270 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_271 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_272 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_273 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_274 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_275 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_276 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_277 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_278 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_279 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_28 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_280 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_281 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_282 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_283 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_284 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_285 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_286 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_287 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_288 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_289 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_29 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_290 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_291 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_292 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_293 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_294 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_295 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_296 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_297 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_298 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_299 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_3 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_30 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_300 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_301 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_302 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_303 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_304 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_305 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_306 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_307 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_308 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_309 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_31 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_310 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_311 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_312 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_313 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_314 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_315 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_316 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_317 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_318 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_319 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_32 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_320 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_321 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_322 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_323 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_324 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_325 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_326 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_327 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_328 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_329 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_33 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_330 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_331 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_332 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_333 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_334 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_335 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_336 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_337 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_338 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_339 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_34 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_340 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_341 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_342 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_343 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_344 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_345 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_346 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_347 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_348 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_349 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_35 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_350 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_351 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_352 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_353 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_354 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_355 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_356 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_357 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_358 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_359 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_36 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_360 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_361 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_362 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_363 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_364 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_365 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_366 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_367 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_368 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_369 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_37 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_370 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_371 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_372 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_373 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_374 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_375 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_376 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_377 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_378 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_379 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_38 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_380 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_381 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_382 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_383 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_384 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_385 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_386 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_387 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_39 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_4 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_40 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_41 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_42 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_43 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_44 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_45 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_46 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_47 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_48 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_49 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_5 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_50 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_51 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_52 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_53 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_54 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_55 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_56 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_57 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_58 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_59 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_6 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_60 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_61 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_62 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_63 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_64 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_65 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_66 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_67 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_68 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_69 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_7 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_70 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_71 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_72 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_73 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_74 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_75 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_76 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_77 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_78 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_79 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_8 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_80 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_81 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_82 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_83 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_84 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_85 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_86 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_87 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_88 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_89 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_9 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_90 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_91 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_92 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_93 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_94 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_95 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_96 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_97 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_98 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__decap_3 PHY_99 (.VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1000 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1001 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1002 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1003 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1004 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1005 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1006 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1007 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1008 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1009 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1010 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1011 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1012 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1013 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1014 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1015 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1016 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1017 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1018 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1019 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1020 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1021 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1022 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1023 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1024 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1025 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1026 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1027 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1028 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1029 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1030 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1031 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1032 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1033 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1034 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1035 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1036 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1037 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1038 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1039 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1040 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1041 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1042 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1043 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1044 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1045 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1046 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1047 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1048 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1049 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1050 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1051 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1052 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1053 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1054 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1055 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1056 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1057 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1058 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1059 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1060 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1061 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1062 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1063 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1064 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1065 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1066 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1067 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1068 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1069 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1070 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1071 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1072 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1073 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1074 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1075 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1076 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1077 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1078 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1079 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1080 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1081 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1082 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1083 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1084 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1085 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1086 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1087 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1088 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1089 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1090 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1091 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1092 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1093 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1094 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1095 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1096 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1097 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1098 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1099 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1100 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1101 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1102 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1103 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1104 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1105 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1106 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1107 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1108 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1109 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1110 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1111 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1112 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1113 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1114 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1115 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1116 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1117 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1118 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1119 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1120 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1121 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1122 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1123 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1124 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1125 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1126 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1127 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1128 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1129 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1130 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1131 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1132 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1133 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1134 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1135 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1136 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1137 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1138 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1139 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1140 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1141 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1142 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1143 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1144 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1145 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1146 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1147 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1148 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1149 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1150 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1151 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1152 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1153 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1154 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1155 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1156 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1157 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1158 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1159 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1160 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1161 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1162 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1163 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1164 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1165 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1166 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1167 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1168 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1169 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1170 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1171 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1172 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1173 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1174 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1175 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1176 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1177 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1178 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1179 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1180 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1181 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1182 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1183 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1184 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1185 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1186 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1187 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1188 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1189 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1190 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1191 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1192 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1193 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1194 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1195 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1196 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1197 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1198 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1199 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1200 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1201 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1202 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1203 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1204 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1205 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1206 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1207 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1208 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1209 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1210 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1211 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1212 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1213 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1214 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1215 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1216 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1217 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1218 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1219 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1220 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1221 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1222 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1223 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1224 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1225 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1226 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1227 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1228 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1229 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1230 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1231 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1232 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1233 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1234 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1235 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1236 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1237 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1238 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1239 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1240 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1241 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1242 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1243 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1244 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1245 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1246 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1247 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1248 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1249 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1250 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1251 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1252 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1253 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1254 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1255 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1256 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1257 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1258 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1259 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1260 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1261 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1262 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1263 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1264 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1265 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1266 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1267 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1268 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1269 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1270 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1271 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1272 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1273 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1274 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1275 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1276 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1277 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1278 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1279 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1280 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1281 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1282 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1283 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1284 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1285 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1286 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1287 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1288 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1289 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1290 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1291 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1292 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1293 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1294 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1295 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1296 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1297 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1298 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1299 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1300 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1301 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1302 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1303 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1304 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1305 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1306 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1307 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1308 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1309 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1310 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1311 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1312 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1313 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1314 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1315 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1316 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1317 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1318 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1319 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1320 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1321 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1322 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1323 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1324 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1325 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1326 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1327 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1328 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1329 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1330 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1331 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1332 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1333 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1334 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1335 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1336 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1337 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1338 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1339 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1340 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1341 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1342 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1343 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1344 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1345 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1346 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1347 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1348 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1349 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1350 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1351 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1352 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1353 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1354 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1355 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1356 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1357 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1358 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1359 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1360 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1361 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1362 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1363 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1364 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1365 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1366 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1367 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1368 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1369 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1370 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1371 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1372 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1373 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1374 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1375 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1376 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1377 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1378 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1379 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1380 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1381 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1382 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1383 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1384 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1385 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1386 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1387 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1388 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1389 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1390 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1391 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1392 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1393 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1394 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1395 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1396 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1397 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1398 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1399 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1400 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1401 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1402 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1403 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1404 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1405 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1406 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1407 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1408 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1409 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1410 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1411 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1412 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1413 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1414 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1415 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1416 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1417 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1418 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1419 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1420 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1421 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1422 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1423 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1424 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1425 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1426 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1427 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1428 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1429 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1430 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1431 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1432 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1433 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1434 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1435 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1436 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1437 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1438 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1439 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1440 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1441 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1442 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1443 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1444 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1445 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1446 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1447 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1448 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1449 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1450 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1451 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1452 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1453 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1454 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1455 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1456 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1457 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1458 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1459 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1460 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1461 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1462 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1463 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1464 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1465 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1466 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1467 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1468 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1469 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1470 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1471 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1472 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1473 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1474 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1475 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1476 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1477 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1478 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1479 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1480 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1481 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1482 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1483 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1484 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1485 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1486 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1487 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1488 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1489 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1490 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1491 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1492 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1493 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1494 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1495 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1496 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1497 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1498 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1499 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1500 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1501 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1502 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1503 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1504 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1505 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1506 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1507 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1508 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1509 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1510 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1511 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1512 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1513 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1514 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1515 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1516 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1517 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1518 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1519 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1520 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1521 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1522 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1523 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1524 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1525 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1526 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1527 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1528 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1529 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1530 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1531 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1532 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1533 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1534 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1535 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1536 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1537 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1538 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1539 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1540 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1541 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1542 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1543 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1544 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1545 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1546 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1547 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1548 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1549 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1550 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1551 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1552 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1553 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1554 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1555 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1556 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1557 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1558 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1559 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1560 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1561 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1562 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1563 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1564 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1565 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1566 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1567 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1568 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1569 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1570 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1571 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1572 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1573 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1574 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1575 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1576 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1577 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1578 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1579 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1580 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1581 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1582 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1583 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1584 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1585 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1586 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1587 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1588 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1589 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1590 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1591 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1592 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1593 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1594 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1595 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1596 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1597 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1598 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1599 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1600 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1601 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1602 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1603 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1604 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1605 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1606 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1607 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1608 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1609 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1610 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1611 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1612 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1613 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1614 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1615 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1616 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1617 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1618 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1619 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1620 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1621 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1622 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1623 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1624 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1625 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1626 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1627 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1628 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1629 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1630 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1631 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1632 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1633 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1634 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1635 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1636 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1637 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1638 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1639 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1640 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1641 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1642 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1643 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1644 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1645 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1646 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1647 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1648 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1649 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1650 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1651 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1652 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1653 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1654 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1655 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1656 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1657 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1658 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1659 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1660 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1661 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1662 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1663 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1664 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1665 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1666 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1667 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1668 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1669 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1670 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1671 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1672 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1673 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1674 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1675 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1676 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1677 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1678 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1679 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1680 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1681 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1682 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1683 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1684 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1685 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1686 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1687 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1688 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1689 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1690 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1691 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1692 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1693 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1694 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1695 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1696 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1697 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1698 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1699 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1700 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1701 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1702 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1703 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1704 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1705 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1706 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1707 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1708 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1709 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1710 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1711 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1712 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1713 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1714 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1715 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1716 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1717 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1718 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1719 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1720 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1721 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1722 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1723 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1724 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1725 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1726 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1727 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1728 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1729 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1730 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1731 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1732 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1733 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1734 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1735 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1736 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1737 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1738 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1739 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1740 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1741 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1742 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1743 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1744 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1745 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1746 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1747 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1748 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1749 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1750 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1751 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1752 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1753 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1754 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1755 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1756 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1757 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1758 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1759 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1760 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1761 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1762 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1763 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1764 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1765 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1766 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1767 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1768 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1769 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1770 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1771 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1772 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1773 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1774 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1775 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1776 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1777 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1778 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1779 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1780 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1781 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1782 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1783 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1784 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1785 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1786 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1787 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1788 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1789 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1790 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1791 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1792 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1793 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1794 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1795 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1796 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1797 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1798 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1799 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1800 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1801 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1802 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1803 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1804 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1805 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1806 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1807 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1808 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1809 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1810 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1811 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1812 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1813 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1814 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1815 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1816 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1817 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1818 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1819 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1820 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1821 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1822 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1823 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1824 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1825 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1826 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1827 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1828 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1829 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1830 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1831 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1832 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1833 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1834 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1835 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1836 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1837 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1838 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1839 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1840 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1841 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1842 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1843 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1844 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1845 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1846 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1847 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1848 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1849 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1850 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1851 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1852 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1853 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1854 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1855 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1856 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1857 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1858 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1859 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1860 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1861 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1862 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1863 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1864 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1865 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1866 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1867 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1868 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1869 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1870 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1871 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1872 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1873 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1874 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1875 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1876 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1877 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1878 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1879 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1880 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1881 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1882 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1883 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1884 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1885 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1886 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1887 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1888 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1889 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1890 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1891 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1892 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1893 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1894 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1895 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1896 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1897 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1898 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1899 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1900 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1901 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1902 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1903 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1904 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1905 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1906 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1907 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1908 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1909 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1910 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1911 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1912 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1913 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1914 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1915 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1916 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1917 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1918 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1919 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1920 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1921 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1922 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1923 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1924 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1925 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1926 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1927 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1928 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1929 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1930 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1931 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1932 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1933 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1934 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1935 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1936 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1937 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1938 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1939 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1940 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1941 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1942 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1943 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1944 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1945 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1946 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1947 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1948 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1949 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1950 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1951 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1952 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1953 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1954 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1955 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1956 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1957 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1958 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1959 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1960 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1961 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1962 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1963 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1964 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1965 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1966 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1967 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1968 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1969 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1970 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1971 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1972 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1973 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1974 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1975 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1976 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1977 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1978 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1979 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1980 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1981 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1982 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1983 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1984 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1985 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1986 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1987 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1988 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1989 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1990 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1991 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1992 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1993 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1994 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1995 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1996 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1997 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1998 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1999 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2000 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2001 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2002 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2003 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2004 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2005 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2006 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2007 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2008 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2009 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2010 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2011 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2012 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2013 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2014 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2015 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2016 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2017 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2018 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2019 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2020 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2021 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2022 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2023 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2024 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2025 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2026 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2027 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2028 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2029 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2030 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2031 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2032 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2033 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2034 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2035 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2036 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2037 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2038 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2039 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2040 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2041 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2042 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2043 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2044 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2045 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2046 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2047 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2048 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2049 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2050 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2051 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2052 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2053 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2054 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2055 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2056 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2057 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2058 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2059 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2060 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2061 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2062 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2063 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2064 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2065 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2066 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2067 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2068 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2069 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2070 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2071 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2072 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2073 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2074 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2075 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2076 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2077 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2078 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2079 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2080 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2081 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2082 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2083 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2084 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2085 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2086 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2087 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2088 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2089 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2090 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2091 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2092 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2093 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2094 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2095 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2096 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2097 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2098 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2099 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2100 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2101 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2102 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2103 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2104 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2105 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2106 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2107 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2108 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2109 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2110 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2111 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2112 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2113 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2114 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2115 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2116 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2117 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2118 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2119 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2120 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2121 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2122 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2123 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2124 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2125 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2126 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2127 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2128 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2129 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2130 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2131 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2132 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2133 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2134 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2135 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2136 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2137 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2138 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2139 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2140 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2141 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2142 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2143 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2144 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2145 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2146 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2147 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2148 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2149 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2150 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2151 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_388 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_389 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_390 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_391 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_392 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_393 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_394 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_395 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_396 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_397 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_398 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_399 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_400 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_401 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_402 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_403 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_404 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_405 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_406 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_407 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_408 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_409 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_410 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_411 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_412 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_413 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_414 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_415 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_416 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_417 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_418 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_419 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_420 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_421 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_422 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_423 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_424 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_425 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_426 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_427 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_428 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_429 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_430 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_431 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_432 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_433 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_434 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_435 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_436 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_437 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_438 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_439 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_440 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_441 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_442 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_443 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_444 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_445 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_446 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_447 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_448 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_449 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_450 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_451 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_452 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_453 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_454 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_455 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_456 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_457 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_458 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_459 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_460 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_461 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_462 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_463 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_464 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_465 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_466 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_467 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_468 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_469 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_470 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_471 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_472 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_473 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_474 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_475 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_476 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_477 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_478 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_479 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_480 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_481 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_482 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_483 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_484 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_485 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_486 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_487 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_488 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_489 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_490 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_491 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_492 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_493 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_494 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_495 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_496 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_497 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_498 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_499 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_500 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_501 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_502 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_503 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_504 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_505 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_506 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_507 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_508 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_509 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_510 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_511 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_512 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_513 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_514 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_515 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_516 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_517 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_518 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_519 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_520 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_521 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_522 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_523 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_524 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_525 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_526 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_527 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_528 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_529 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_530 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_531 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_532 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_533 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_534 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_535 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_536 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_537 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_538 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_539 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_540 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_541 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_542 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_543 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_544 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_545 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_546 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_547 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_548 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_549 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_550 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_551 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_552 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_553 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_554 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_555 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_556 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_557 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_558 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_559 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_560 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_561 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_562 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_563 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_564 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_565 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_566 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_567 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_568 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_569 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_570 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_571 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_572 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_573 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_574 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_575 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_576 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_577 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_578 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_579 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_580 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_581 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_582 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_583 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_584 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_585 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_586 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_587 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_588 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_589 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_590 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_591 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_592 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_593 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_594 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_595 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_596 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_597 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_598 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_599 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_600 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_601 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_602 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_603 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_604 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_605 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_606 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_607 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_608 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_609 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_610 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_611 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_612 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_613 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_614 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_615 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_616 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_617 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_618 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_619 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_620 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_621 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_622 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_623 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_624 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_625 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_626 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_627 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_628 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_629 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_630 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_631 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_632 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_633 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_634 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_635 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_636 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_637 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_638 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_639 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_640 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_641 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_642 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_643 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_644 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_645 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_646 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_647 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_648 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_649 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_650 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_651 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_652 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_653 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_654 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_655 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_656 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_657 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_658 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_659 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_660 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_661 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_662 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_663 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_664 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_665 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_666 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_667 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_668 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_669 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_670 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_671 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_672 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_673 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_674 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_675 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_676 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_677 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_678 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_679 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_680 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_681 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_682 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_683 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_684 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_685 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_686 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_687 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_688 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_689 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_690 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_691 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_692 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_693 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_694 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_695 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_696 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_697 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_698 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_699 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_700 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_701 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_702 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_703 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_704 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_705 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_706 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_707 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_708 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_709 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_710 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_711 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_712 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_713 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_714 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_715 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_716 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_717 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_718 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_719 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_720 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_721 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_722 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_723 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_724 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_725 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_726 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_727 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_728 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_729 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_730 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_731 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_732 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_733 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_734 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_735 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_736 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_737 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_738 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_739 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_740 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_741 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_742 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_743 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_744 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_745 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_746 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_747 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_748 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_749 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_750 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_751 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_752 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_753 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_754 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_755 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_756 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_757 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_758 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_759 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_760 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_761 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_762 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_763 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_764 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_765 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_766 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_767 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_768 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_769 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_770 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_771 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_772 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_773 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_774 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_775 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_776 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_777 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_778 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_779 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_780 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_781 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_782 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_783 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_784 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_785 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_786 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_787 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_788 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_789 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_790 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_791 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_792 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_793 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_794 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_795 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_796 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_797 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_798 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_799 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_800 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_801 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_802 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_803 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_804 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_805 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_806 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_807 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_808 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_809 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_810 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_811 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_812 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_813 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_814 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_815 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_816 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_817 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_818 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_819 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_820 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_821 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_822 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_823 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_824 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_825 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_826 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_827 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_828 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_829 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_830 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_831 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_832 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_833 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_834 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_835 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_836 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_837 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_838 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_839 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_840 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_841 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_842 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_843 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_844 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_845 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_846 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_847 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_848 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_849 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_850 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_851 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_852 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_853 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_854 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_855 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_856 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_857 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_858 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_859 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_860 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_861 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_862 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_863 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_864 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_865 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_866 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_867 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_868 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_869 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_870 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_871 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_872 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_873 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_874 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_875 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_876 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_877 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_878 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_879 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_880 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_881 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_882 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_883 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_884 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_885 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_886 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_887 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_888 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_889 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_890 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_891 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_892 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_893 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_894 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_895 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_896 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_897 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_898 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_899 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_900 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_901 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_902 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_903 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_904 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_905 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_906 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_907 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_908 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_909 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_910 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_911 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_912 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_913 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_914 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_915 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_916 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_917 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_918 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_919 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_920 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_921 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_922 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_923 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_924 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_925 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_926 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_927 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_928 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_929 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_930 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_931 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_932 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_933 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_934 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_935 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_936 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_937 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_938 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_939 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_940 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_941 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_942 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_943 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_944 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_945 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_946 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_947 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_948 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_949 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_950 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_951 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_952 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_953 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_954 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_955 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_956 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_957 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_958 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_959 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_960 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_961 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_962 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_963 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_964 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_965 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_966 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_967 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_968 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_969 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_970 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_971 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_972 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_973 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_974 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_975 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_976 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_977 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_978 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_979 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_980 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_981 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_982 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_983 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_984 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_985 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_986 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_987 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_988 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_989 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_990 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_991 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_992 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_993 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_994 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_995 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_996 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_997 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_998 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_999 (.VGND(vssa1),
    .VPWR(vdda1));
 sky130_fd_sc_hd__dfxtp_2 _0_ (.CLK(clknet_1_1__leaf_Vref),
    .D(DIn1[7]),
    .VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1),
    .Q(Vout2));
 sky130_fd_sc_hd__dfxtp_2 _1_ (.CLK(clknet_1_1__leaf_Vref),
    .D(DIn2[7]),
    .VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1),
    .Q(Vout3));
 sky130_fd_sc_hd__dfxtp_2 _2_ (.CLK(clknet_1_0__leaf_Vref),
    .D(DIn0[0]),
    .VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1),
    .Q(Vout0));
 sky130_fd_sc_hd__dfxtp_2 _3_ (.CLK(clknet_1_0__leaf_Vref),
    .D(DIn1[0]),
    .VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1),
    .Q(Vout1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_Vref (.A(Vref),
    .VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1),
    .X(clknet_0_Vref));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_Vref (.A(clknet_0_Vref),
    .VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1),
    .X(clknet_1_0__leaf_Vref));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_Vref (.A(clknet_0_Vref),
    .VGND(vssa1),
    .VNB(vssa1),
    .VPB(vdda1),
    .VPWR(vdda1),
    .X(clknet_1_1__leaf_Vref));
endmodule
