* /home/dinesha/workarea/opencore/git/8bit_dac/schematics/switch/switch.cir


.lib "../sky130_fd_pr/models/sky130.lib.spice" tt

xM3  Net-_M3-Pad1_ Net-_M1-Pad1_ vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5		
xM4  Net-_M3-Pad1_ Net-_M1-Pad1_ GND GND sky130_fd_pr__nfet_01v8 w=0.42 l=0.5		
xM1  Net-_M1-Pad1_ digital_input vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5		
xM2  Net-_M1-Pad1_ digital_input GND GND sky130_fd_pr__nfet_01v8 w=0.42 l=0.5		
xM6  Vout Net-_M1-Pad1_ vin_2 GND sky130_fd_pr__nfet_01v8 w=0.42 l=0.5		
xM5  Vout Net-_M1-Pad1_ vin_1 vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5		
xM7  vin_1 Net-_M3-Pad1_ Vout GND sky130_fd_pr__nfet_01v8 w=0.42 l=0.5		
xM8  vin_2 Net-_M3-Pad1_ Vout vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5		


Vdd vdd 0 3.3
Vin_1 vin_1 0 2.5
Vin_2 vin_2 0 2
Vd0 digital_input 0 pulse (0 1.8 0s 0s 0s 5us 10us)

.tran 0.1us 40us

.control
run

plot V(vin_1) V(vin_2) V(digital_input) V(vout)

.endc



.end
