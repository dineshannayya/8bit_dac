* C:\FOSSEE\eSim\library\SubcircuitLibrary\switch\switch.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 04/19/23 16:38:01

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
M6  Net-_M5-Pad1_ Net-_M1-Pad1_ /vdd /vdd mosfet_p		
M5  Net-_M5-Pad1_ Net-_M1-Pad1_ GND GND mosfet_n		
M2  Net-_M1-Pad1_ /digital_input /vdd /vdd mosfet_p		
M1  Net-_M1-Pad1_ /digital_input GND GND mosfet_n		
M3  /Vout Net-_M1-Pad1_ /vrefl GND mosfet_n		
M4  /Vout Net-_M1-Pad1_ /vrefh /vdd mosfet_p		
M8  /vrefh Net-_M5-Pad1_ /Vout GND mosfet_n		
M7  /vrefl Net-_M5-Pad1_ /Vout /vdd mosfet_p		
U1  /vdd /digital_input /vrefh /vrefl /Vout PORT		

.end
