* D:\vlsi\github\8bit_dac\schematics\2bit_DAC\2bit_DAC.cir

.include switch.sub

.subckt resistor b a VSUBS
X0 a b VSUBS sky130_fd_pr__res_generic_nd w=160000u l=820000u
.ends

xR4  Net-_R3-Pad2_ vrefl VSUBS resistor
xR3  Net-_R2-Pad2_ Net-_R3-Pad2_ VSUBS resistor
xR2  Net-_R1-Pad2_ Net-_R2-Pad2_ VSUBS resistor
xR1  vrefh Net-_R1-Pad2_ VSUBS resistor
xS2  vdd d0 Net-_R3-Pad2_ vrefl Net1 switch		
xS1  vdd d0 Net-_R1-Pad2_ Net-_R2-Pad2_ Net2 switch		
xS3  vdd d1 Net1 Net2 vout switch		

Vdd vdd 0 3.3
Vrefh vrefh 0 3.3
Vrefl vrefl 0 0.0
Vd0 d0 0 pulse(0 1.8 0ns 0.1ns 0.1ns 5us 10us)
Vd1 d1 0 pulse(0 1.8 0ns 0.1ns 0.1ns 10us 20us)

.tran 0.1us 80us

.control
run

plot V(d0) V(d1) v(vout)

.endc

.end
